//Generated from netlist by SpyDrNet
//netlist name: SDN_VERILOG_NETLIST_logical_tile_io_mode_physical__iopad
module fpga_top
(
    reset,
    clk,
    gfpga_pad_GPIO_PAD,
    bl,
    wl
);

    input reset;
    input clk;
    inout [0:127]gfpga_pad_GPIO_PAD;
    input [0:21507]bl;
    input [0:21507]wl;

    wire reset;
    wire clk;
    wire [0:127]gfpga_pad_GPIO_PAD;
    wire [0:21507]bl;
    wire [0:21507]wl;
    wire [0:19]cbx_1__0__0_chanx_left_out;
    wire [0:19]cbx_1__0__0_chanx_right_out;
    wire [0:19]cbx_1__0__1_chanx_left_out;
    wire [0:19]cbx_1__0__1_chanx_right_out;
    wire [0:19]cbx_1__0__2_chanx_left_out;
    wire [0:19]cbx_1__0__2_chanx_right_out;
    wire [0:19]cbx_1__0__3_chanx_left_out;
    wire [0:19]cbx_1__0__3_chanx_right_out;
    wire [0:19]cbx_1__1__0_chanx_left_out;
    wire [0:19]cbx_1__1__0_chanx_right_out;
    wire [0:19]cbx_1__1__10_chanx_left_out;
    wire [0:19]cbx_1__1__10_chanx_right_out;
    wire [0:19]cbx_1__1__11_chanx_left_out;
    wire [0:19]cbx_1__1__11_chanx_right_out;
    wire [0:19]cbx_1__1__1_chanx_left_out;
    wire [0:19]cbx_1__1__1_chanx_right_out;
    wire [0:19]cbx_1__1__2_chanx_left_out;
    wire [0:19]cbx_1__1__2_chanx_right_out;
    wire [0:19]cbx_1__1__3_chanx_left_out;
    wire [0:19]cbx_1__1__3_chanx_right_out;
    wire [0:19]cbx_1__1__4_chanx_left_out;
    wire [0:19]cbx_1__1__4_chanx_right_out;
    wire [0:19]cbx_1__1__5_chanx_left_out;
    wire [0:19]cbx_1__1__5_chanx_right_out;
    wire [0:19]cbx_1__1__6_chanx_left_out;
    wire [0:19]cbx_1__1__6_chanx_right_out;
    wire [0:19]cbx_1__1__7_chanx_left_out;
    wire [0:19]cbx_1__1__7_chanx_right_out;
    wire [0:19]cbx_1__1__8_chanx_left_out;
    wire [0:19]cbx_1__1__8_chanx_right_out;
    wire [0:19]cbx_1__1__9_chanx_left_out;
    wire [0:19]cbx_1__1__9_chanx_right_out;
    wire [0:19]cbx_1__4__0_chanx_left_out;
    wire [0:19]cbx_1__4__0_chanx_right_out;
    wire [0:19]cbx_1__4__1_chanx_left_out;
    wire [0:19]cbx_1__4__1_chanx_right_out;
    wire [0:19]cbx_1__4__2_chanx_left_out;
    wire [0:19]cbx_1__4__2_chanx_right_out;
    wire [0:19]cbx_1__4__3_chanx_left_out;
    wire [0:19]cbx_1__4__3_chanx_right_out;
    wire [0:19]cby_0__1__0_chany_bottom_out;
    wire [0:19]cby_0__1__0_chany_top_out;
    wire [0:19]cby_0__1__1_chany_bottom_out;
    wire [0:19]cby_0__1__1_chany_top_out;
    wire [0:19]cby_0__1__2_chany_bottom_out;
    wire [0:19]cby_0__1__2_chany_top_out;
    wire [0:19]cby_0__1__3_chany_bottom_out;
    wire [0:19]cby_0__1__3_chany_top_out;
    wire [0:19]cby_1__1__0_chany_bottom_out;
    wire [0:19]cby_1__1__0_chany_top_out;
    wire [0:19]cby_1__1__10_chany_bottom_out;
    wire [0:19]cby_1__1__10_chany_top_out;
    wire [0:19]cby_1__1__11_chany_bottom_out;
    wire [0:19]cby_1__1__11_chany_top_out;
    wire [0:19]cby_1__1__1_chany_bottom_out;
    wire [0:19]cby_1__1__1_chany_top_out;
    wire [0:19]cby_1__1__2_chany_bottom_out;
    wire [0:19]cby_1__1__2_chany_top_out;
    wire [0:19]cby_1__1__3_chany_bottom_out;
    wire [0:19]cby_1__1__3_chany_top_out;
    wire [0:19]cby_1__1__4_chany_bottom_out;
    wire [0:19]cby_1__1__4_chany_top_out;
    wire [0:19]cby_1__1__5_chany_bottom_out;
    wire [0:19]cby_1__1__5_chany_top_out;
    wire [0:19]cby_1__1__6_chany_bottom_out;
    wire [0:19]cby_1__1__6_chany_top_out;
    wire [0:19]cby_1__1__7_chany_bottom_out;
    wire [0:19]cby_1__1__7_chany_top_out;
    wire [0:19]cby_1__1__8_chany_bottom_out;
    wire [0:19]cby_1__1__8_chany_top_out;
    wire [0:19]cby_1__1__9_chany_bottom_out;
    wire [0:19]cby_1__1__9_chany_top_out;
    wire [0:19]cby_4__1__0_chany_bottom_out;
    wire [0:19]cby_4__1__0_chany_top_out;
    wire [0:19]cby_4__1__1_chany_bottom_out;
    wire [0:19]cby_4__1__1_chany_top_out;
    wire [0:19]cby_4__1__2_chany_bottom_out;
    wire [0:19]cby_4__1__2_chany_top_out;
    wire [0:19]cby_4__1__3_chany_bottom_out;
    wire [0:19]cby_4__1__3_chany_top_out;
    wire [0:19]sb_0__0__0_chanx_right_out;
    wire [0:19]sb_0__0__0_chany_top_out;
    wire [0:19]sb_0__1__0_chanx_right_out;
    wire [0:19]sb_0__1__0_chany_bottom_out;
    wire [0:19]sb_0__1__0_chany_top_out;
    wire [0:19]sb_0__1__1_chanx_right_out;
    wire [0:19]sb_0__1__1_chany_bottom_out;
    wire [0:19]sb_0__1__1_chany_top_out;
    wire [0:19]sb_0__1__2_chanx_right_out;
    wire [0:19]sb_0__1__2_chany_bottom_out;
    wire [0:19]sb_0__1__2_chany_top_out;
    wire [0:19]sb_0__4__0_chanx_right_out;
    wire [0:19]sb_0__4__0_chany_bottom_out;
    wire [0:19]sb_1__0__0_chanx_left_out;
    wire [0:19]sb_1__0__0_chanx_right_out;
    wire [0:19]sb_1__0__0_chany_top_out;
    wire [0:19]sb_1__0__1_chanx_left_out;
    wire [0:19]sb_1__0__1_chanx_right_out;
    wire [0:19]sb_1__0__1_chany_top_out;
    wire [0:19]sb_1__0__2_chanx_left_out;
    wire [0:19]sb_1__0__2_chanx_right_out;
    wire [0:19]sb_1__0__2_chany_top_out;
    wire [0:19]sb_1__1__0_chanx_left_out;
    wire [0:19]sb_1__1__0_chanx_right_out;
    wire [0:19]sb_1__1__0_chany_bottom_out;
    wire [0:19]sb_1__1__0_chany_top_out;
    wire [0:19]sb_1__1__1_chanx_left_out;
    wire [0:19]sb_1__1__1_chanx_right_out;
    wire [0:19]sb_1__1__1_chany_bottom_out;
    wire [0:19]sb_1__1__1_chany_top_out;
    wire [0:19]sb_1__1__2_chanx_left_out;
    wire [0:19]sb_1__1__2_chanx_right_out;
    wire [0:19]sb_1__1__2_chany_bottom_out;
    wire [0:19]sb_1__1__2_chany_top_out;
    wire [0:19]sb_1__1__3_chanx_left_out;
    wire [0:19]sb_1__1__3_chanx_right_out;
    wire [0:19]sb_1__1__3_chany_bottom_out;
    wire [0:19]sb_1__1__3_chany_top_out;
    wire [0:19]sb_1__1__4_chanx_left_out;
    wire [0:19]sb_1__1__4_chanx_right_out;
    wire [0:19]sb_1__1__4_chany_bottom_out;
    wire [0:19]sb_1__1__4_chany_top_out;
    wire [0:19]sb_1__1__5_chanx_left_out;
    wire [0:19]sb_1__1__5_chanx_right_out;
    wire [0:19]sb_1__1__5_chany_bottom_out;
    wire [0:19]sb_1__1__5_chany_top_out;
    wire [0:19]sb_1__1__6_chanx_left_out;
    wire [0:19]sb_1__1__6_chanx_right_out;
    wire [0:19]sb_1__1__6_chany_bottom_out;
    wire [0:19]sb_1__1__6_chany_top_out;
    wire [0:19]sb_1__1__7_chanx_left_out;
    wire [0:19]sb_1__1__7_chanx_right_out;
    wire [0:19]sb_1__1__7_chany_bottom_out;
    wire [0:19]sb_1__1__7_chany_top_out;
    wire [0:19]sb_1__1__8_chanx_left_out;
    wire [0:19]sb_1__1__8_chanx_right_out;
    wire [0:19]sb_1__1__8_chany_bottom_out;
    wire [0:19]sb_1__1__8_chany_top_out;
    wire [0:19]sb_1__4__0_chanx_left_out;
    wire [0:19]sb_1__4__0_chanx_right_out;
    wire [0:19]sb_1__4__0_chany_bottom_out;
    wire [0:19]sb_1__4__1_chanx_left_out;
    wire [0:19]sb_1__4__1_chanx_right_out;
    wire [0:19]sb_1__4__1_chany_bottom_out;
    wire [0:19]sb_1__4__2_chanx_left_out;
    wire [0:19]sb_1__4__2_chanx_right_out;
    wire [0:19]sb_1__4__2_chany_bottom_out;
    wire [0:19]sb_4__0__0_chanx_left_out;
    wire [0:19]sb_4__0__0_chany_top_out;
    wire [0:19]sb_4__1__0_chanx_left_out;
    wire [0:19]sb_4__1__0_chany_bottom_out;
    wire [0:19]sb_4__1__0_chany_top_out;
    wire [0:19]sb_4__1__1_chanx_left_out;
    wire [0:19]sb_4__1__1_chany_bottom_out;
    wire [0:19]sb_4__1__1_chany_top_out;
    wire [0:19]sb_4__1__2_chanx_left_out;
    wire [0:19]sb_4__1__2_chany_bottom_out;
    wire [0:19]sb_4__1__2_chany_top_out;
    wire [0:19]sb_4__4__0_chanx_left_out;
    wire [0:19]sb_4__4__0_chany_bottom_out;
    wire [0:9]grid_clb_1__1__grid_left_in;
    wire [0:9]grid_clb_1__1__grid_top_in;
    wire [0:9]grid_clb_1__1__grid_right_in;
    wire [0:9]grid_clb_1__1__grid_bottom_in;
    wire [0:9]grid_clb_1__2__grid_left_in;
    wire [0:9]grid_clb_1__2__grid_top_in;
    wire [0:9]grid_clb_1__2__grid_right_in;
    wire [0:9]grid_clb_1__2__grid_bottom_in;
    wire [0:9]grid_clb_1__3__grid_left_in;
    wire [0:9]grid_clb_1__3__grid_top_in;
    wire [0:9]grid_clb_1__3__grid_right_in;
    wire [0:9]grid_clb_1__3__grid_bottom_in;
    wire [0:9]grid_clb_1__4__grid_left_in;
    wire [0:9]grid_clb_1__4__grid_top_in;
    wire [0:9]grid_clb_1__4__grid_right_in;
    wire [0:9]grid_clb_1__4__grid_bottom_in;
    wire [0:9]grid_clb_2__1__grid_left_in;
    wire [0:9]grid_clb_2__1__grid_top_in;
    wire [0:9]grid_clb_2__1__grid_right_in;
    wire [0:9]grid_clb_2__1__grid_bottom_in;
    wire [0:9]grid_clb_2__2__grid_left_in;
    wire [0:9]grid_clb_2__2__grid_top_in;
    wire [0:9]grid_clb_2__2__grid_right_in;
    wire [0:9]grid_clb_2__2__grid_bottom_in;
    wire [0:9]grid_clb_2__3__grid_left_in;
    wire [0:9]grid_clb_2__3__grid_top_in;
    wire [0:9]grid_clb_2__3__grid_right_in;
    wire [0:9]grid_clb_2__3__grid_bottom_in;
    wire [0:9]grid_clb_2__4__grid_left_in;
    wire [0:9]grid_clb_2__4__grid_top_in;
    wire [0:9]grid_clb_2__4__grid_right_in;
    wire [0:9]grid_clb_2__4__grid_bottom_in;
    wire [0:9]grid_clb_3__1__grid_left_in;
    wire [0:9]grid_clb_3__1__grid_top_in;
    wire [0:9]grid_clb_3__1__grid_right_in;
    wire [0:9]grid_clb_3__1__grid_bottom_in;
    wire [0:9]grid_clb_3__2__grid_left_in;
    wire [0:9]grid_clb_3__2__grid_top_in;
    wire [0:9]grid_clb_3__2__grid_right_in;
    wire [0:9]grid_clb_3__2__grid_bottom_in;
    wire [0:9]grid_clb_3__3__grid_left_in;
    wire [0:9]grid_clb_3__3__grid_top_in;
    wire [0:9]grid_clb_3__3__grid_right_in;
    wire [0:9]grid_clb_3__3__grid_bottom_in;
    wire [0:9]grid_clb_3__4__grid_left_in;
    wire [0:9]grid_clb_3__4__grid_top_in;
    wire [0:9]grid_clb_3__4__grid_right_in;
    wire [0:9]grid_clb_3__4__grid_bottom_in;
    wire [0:9]grid_clb_4__1__grid_left_in;
    wire [0:9]grid_clb_4__1__grid_top_in;
    wire [0:9]grid_clb_4__1__grid_right_in;
    wire [0:9]grid_clb_4__1__grid_bottom_in;
    wire [0:9]grid_clb_4__2__grid_left_in;
    wire [0:9]grid_clb_4__2__grid_top_in;
    wire [0:9]grid_clb_4__2__grid_right_in;
    wire [0:9]grid_clb_4__2__grid_bottom_in;
    wire [0:9]grid_clb_4__3__grid_left_in;
    wire [0:9]grid_clb_4__3__grid_top_in;
    wire [0:9]grid_clb_4__3__grid_right_in;
    wire [0:9]grid_clb_4__3__grid_bottom_in;
    wire [0:9]grid_clb_4__4__grid_left_in;
    wire [0:9]grid_clb_4__4__grid_top_in;
    wire [0:9]grid_clb_4__4__grid_right_in;
    wire [0:9]grid_clb_4__4__grid_bottom_in;
    wire [0:7]grid_io_top_1__5__io_bottom_in;
    wire [0:7]grid_io_top_1__5__io_bottom_out;
    wire [0:7]grid_io_top_2__5__io_bottom_in;
    wire [0:7]grid_io_top_2__5__io_bottom_out;
    wire [0:7]grid_io_top_3__5__io_bottom_in;
    wire [0:7]grid_io_top_3__5__io_bottom_out;
    wire [0:7]grid_io_top_4__5__io_bottom_in;
    wire [0:7]grid_io_top_4__5__io_bottom_out;
    wire [0:7]grid_io_right_5__4__io_left_in;
    wire [0:7]grid_io_right_5__4__io_left_out;
    wire [0:7]grid_io_right_5__3__io_left_in;
    wire [0:7]grid_io_right_5__3__io_left_out;
    wire [0:7]grid_io_right_5__2__io_left_in;
    wire [0:7]grid_io_right_5__2__io_left_out;
    wire [0:7]grid_io_right_5__1__io_left_in;
    wire [0:7]grid_io_right_5__1__io_left_out;
    wire [0:7]grid_io_bottom_4__0__io_top_in;
    wire [0:7]grid_io_bottom_4__0__io_top_out;
    wire [0:7]grid_io_bottom_3__0__io_top_in;
    wire [0:7]grid_io_bottom_3__0__io_top_out;
    wire [0:7]grid_io_bottom_2__0__io_top_in;
    wire [0:7]grid_io_bottom_2__0__io_top_out;
    wire [0:7]grid_io_bottom_1__0__io_top_in;
    wire [0:7]grid_io_bottom_1__0__io_top_out;
    wire [0:7]grid_io_left_0__1__io_right_in;
    wire [0:7]grid_io_left_0__1__io_right_out;
    wire [0:7]grid_io_left_0__2__io_right_in;
    wire [0:7]grid_io_left_0__2__io_right_out;
    wire [0:7]grid_io_left_0__3__io_right_in;
    wire [0:7]grid_io_left_0__3__io_right_out;
    wire [0:7]grid_io_left_0__4__io_right_in;
    wire [0:7]grid_io_left_0__4__io_right_out;
    wire [0:1]sb_0__0__grid_top_r_in;
    wire [0:1]sb_0__0__grid_right_t_in;
    wire [0:1]sb_0__1__grid_top_r_in;
    wire [0:1]sb_0__1__grid_right_t_in;
    wire [0:2]sb_0__1__grid_right_b_in;
    wire [0:1]sb_0__2__grid_top_r_in;
    wire [0:1]sb_0__2__grid_right_t_in;
    wire [0:2]sb_0__2__grid_right_b_in;
    wire [0:1]sb_0__3__grid_top_r_in;
    wire [0:1]sb_0__3__grid_right_t_in;
    wire [0:2]sb_0__3__grid_right_b_in;
    wire [0:2]sb_0__4__grid_right_b_in;
    wire [0:1]sb_1__0__grid_top_r_in;
    wire [0:2]sb_1__0__grid_top_l_in;
    wire [0:1]sb_1__0__grid_right_t_in;
    wire [0:1]sb_2__0__grid_top_r_in;
    wire [0:2]sb_2__0__grid_top_l_in;
    wire [0:1]sb_2__0__grid_right_t_in;
    wire [0:1]sb_3__0__grid_top_r_in;
    wire [0:2]sb_3__0__grid_top_l_in;
    wire [0:1]sb_3__0__grid_right_t_in;
    wire [0:1]sb_1__1__grid_top_r_in;
    wire [0:2]sb_1__1__grid_top_l_in;
    wire [0:1]sb_1__1__grid_right_t_in;
    wire [0:2]sb_1__1__grid_right_b_in;
    wire [0:1]sb_1__2__grid_top_r_in;
    wire [0:2]sb_1__2__grid_top_l_in;
    wire [0:1]sb_1__2__grid_right_t_in;
    wire [0:2]sb_1__2__grid_right_b_in;
    wire [0:1]sb_1__3__grid_top_r_in;
    wire [0:2]sb_1__3__grid_top_l_in;
    wire [0:1]sb_1__3__grid_right_t_in;
    wire [0:2]sb_1__3__grid_right_b_in;
    wire [0:1]sb_2__1__grid_top_r_in;
    wire [0:2]sb_2__1__grid_top_l_in;
    wire [0:1]sb_2__1__grid_right_t_in;
    wire [0:2]sb_2__1__grid_right_b_in;
    wire [0:1]sb_2__2__grid_top_r_in;
    wire [0:2]sb_2__2__grid_top_l_in;
    wire [0:1]sb_2__2__grid_right_t_in;
    wire [0:2]sb_2__2__grid_right_b_in;
    wire [0:1]sb_2__3__grid_top_r_in;
    wire [0:2]sb_2__3__grid_top_l_in;
    wire [0:1]sb_2__3__grid_right_t_in;
    wire [0:2]sb_2__3__grid_right_b_in;
    wire [0:1]sb_3__1__grid_top_r_in;
    wire [0:2]sb_3__1__grid_top_l_in;
    wire [0:1]sb_3__1__grid_right_t_in;
    wire [0:2]sb_3__1__grid_right_b_in;
    wire [0:1]sb_3__2__grid_top_r_in;
    wire [0:2]sb_3__2__grid_top_l_in;
    wire [0:1]sb_3__2__grid_right_t_in;
    wire [0:2]sb_3__2__grid_right_b_in;
    wire [0:1]sb_3__3__grid_top_r_in;
    wire [0:2]sb_3__3__grid_top_l_in;
    wire [0:1]sb_3__3__grid_right_t_in;
    wire [0:2]sb_3__3__grid_right_b_in;
    wire [0:2]sb_1__4__grid_right_b_in;
    wire [0:2]sb_2__4__grid_right_b_in;
    wire [0:2]sb_3__4__grid_right_b_in;
    wire [0:2]sb_4__0__grid_top_l_in;
    wire [0:2]sb_4__1__grid_top_l_in;
    wire [0:2]sb_4__2__grid_top_l_in;
    wire [0:2]sb_4__3__grid_top_l_in;

    tile tile_2__2_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_0__1__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_0__1__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_0__1__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_1__0__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_1__0__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_1__0__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_0__0__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_0__0__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_0__0__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_0__0__grid_top_r_in[1]),
        .grid_left_in(grid_clb_1__1__grid_left_in),
        .grid_bottom_in(grid_clb_1__1__grid_bottom_in),
        .chanx_left_in(sb_0__1__0_chanx_right_out),
        .chanx_left_out(cbx_1__1__0_chanx_left_out),
        .grid_top_out(grid_clb_1__2__grid_bottom_in),
        .chany_bottom_in(sb_1__0__0_chany_top_out),
        .chany_bottom_out(cby_1__1__0_chany_bottom_out),
        .grid_right_out(grid_clb_2__1__grid_left_in),
        .chany_top_in_0(cby_1__1__1_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__3_chanx_left_out),
        .chany_top_out_0(sb_1__1__0_chany_top_out),
        .chanx_right_out_0(sb_1__1__0_chanx_right_out),
        .grid_top_r_in(sb_1__1__grid_top_r_in),
        .grid_top_l_in(sb_1__1__grid_top_l_in),
        .grid_right_t_in(sb_1__1__grid_right_t_in),
        .grid_right_b_in(sb_1__1__grid_right_b_in),
        .grid_bottom_r_in(sb_1__0__grid_top_r_in),
        .grid_bottom_l_in(sb_1__0__grid_top_l_in),
        .grid_left_t_in(sb_0__1__grid_right_t_in),
        .grid_left_b_in(sb_0__1__grid_right_b_in),
        .bl({bl[1648], bl[1649], bl[1650], bl[1651], bl[1652], bl[1653], bl[1654], bl[1655], bl[1656], bl[1657], bl[1658], bl[1659], bl[1660], bl[1661], bl[1662], bl[1663], bl[1664], bl[1665], bl[1666], bl[1667], bl[1668], bl[1669], bl[1670], bl[1671], bl[1672], bl[1673], bl[1674], bl[1675], bl[1676], bl[1677], bl[1678], bl[1679], bl[1680], bl[1681], bl[1682], bl[1683], bl[1684], bl[1685], bl[1686], bl[1687], bl[1688], bl[1689], bl[1690], bl[1691], bl[1692], bl[1693], bl[1694], bl[1695], bl[1696], bl[1697], bl[1698], bl[1699], bl[1700], bl[1701], bl[1702], bl[1703], bl[1704], bl[1705], bl[1706], bl[1707], bl[1708], bl[1709], bl[1710], bl[1711], bl[1712], bl[1713], bl[1714], bl[1715], bl[1716], bl[1717], bl[1718], bl[1719], bl[1720], bl[1721], bl[1722], bl[1723], bl[1724], bl[1725], bl[1726], bl[1727], bl[1728], bl[1729], bl[1730], bl[1731], bl[1732], bl[1733], bl[1734], bl[1735], bl[1736], bl[1737], bl[1738], bl[1739], bl[1740], bl[1741], bl[1742], bl[1743], bl[1744], bl[1745], bl[1746], bl[1747], bl[1748], bl[1749], bl[1750], bl[1751], bl[1752], bl[1753], bl[1754], bl[1755], bl[1756], bl[1757], bl[1758], bl[1759], bl[1760], bl[1761], bl[1762], bl[1763], bl[1764], bl[1765], bl[1766], bl[1767], bl[1768], bl[1769], bl[1770], bl[1771], bl[1772], bl[1773], bl[1774], bl[1775], bl[1776], bl[1777], bl[1778], bl[1779], bl[1780], bl[1781], bl[1782], bl[1783], bl[1784], bl[1785], bl[1786], bl[1787], bl[1788], bl[1789], bl[1790], bl[1791], bl[1792], bl[1793], bl[1794], bl[1795], bl[1796], bl[1797], bl[1798], bl[1799], bl[1800], bl[1801], bl[1802], bl[1803], bl[1804], bl[1805], bl[1806], bl[1807], bl[1808], bl[1809], bl[1810], bl[1811], bl[1812], bl[1813], bl[1814], bl[1815], bl[1816], bl[1817], bl[1818], bl[1819], bl[1820], bl[1821], bl[1822], bl[1823], bl[1824], bl[1825], bl[1826], bl[1827], bl[1828], bl[1829], bl[1830], bl[1831], bl[1832], bl[1833], bl[1834], bl[1835], bl[1836], bl[1837], bl[1838], bl[1839], bl[1840], bl[1841], bl[1842], bl[1843], bl[1844], bl[1845], bl[1846], bl[1847], bl[1848], bl[1849], bl[1850], bl[1851], bl[1852], bl[1853], bl[1854], bl[1855], bl[1856], bl[1857], bl[1858], bl[1859], bl[1860], bl[1861], bl[1862], bl[1863], bl[1864], bl[1865], bl[1866], bl[1867], bl[1868], bl[1869], bl[1870], bl[1871], bl[1872], bl[1873], bl[1874], bl[1875], bl[1876], bl[1877], bl[1878], bl[1879], bl[1880], bl[1881], bl[1882], bl[1883], bl[1884], bl[1885], bl[1886], bl[1887], bl[1888], bl[1889], bl[1890], bl[1891], bl[1892], bl[1893], bl[1894], bl[1895], bl[1896], bl[1897], bl[1898], bl[1899], bl[1900], bl[1901], bl[1902], bl[1903], bl[1904], bl[1905], bl[1906], bl[1907], bl[1908], bl[1909], bl[1910], bl[1911], bl[1912], bl[1913], bl[1914], bl[1915], bl[1916], bl[1917], bl[1918], bl[1919], bl[1920], bl[1921], bl[1922], bl[1923], bl[1924], bl[1925], bl[1926], bl[1927], bl[1928], bl[1929], bl[1930], bl[1931], bl[1932], bl[1933], bl[1934], bl[1935], bl[1936], bl[1937], bl[1938], bl[1939], bl[1940], bl[1941], bl[1942], bl[1943], bl[1944], bl[1945], bl[1946], bl[1947], bl[1948], bl[1949], bl[1950], bl[1951], bl[1952], bl[1953], bl[1954], bl[1955], bl[1956], bl[1957], bl[1958], bl[1959], bl[1960], bl[1961], bl[1962], bl[1963], bl[1964], bl[1965], bl[1966], bl[1967], bl[1968], bl[1969], bl[1970], bl[1971], bl[1972], bl[1973], bl[1974], bl[1975], bl[1976], bl[1977], bl[1978], bl[1979], bl[1980], bl[1981], bl[1982], bl[1983], bl[1984], bl[1985], bl[1986], bl[1987], bl[1988], bl[1989], bl[1990], bl[1991], bl[1992], bl[1993], bl[1994], bl[1995], bl[1996], bl[1997], bl[1998], bl[1999], bl[2000], bl[2001], bl[2002], bl[2003], bl[2004], bl[2005], bl[2006], bl[2007], bl[2008], bl[2009], bl[2010], bl[2011], bl[2012], bl[2013], bl[2014], bl[2015], bl[2016], bl[2017], bl[2018], bl[2019], bl[2020], bl[2021], bl[2022], bl[2023], bl[2024], bl[2025], bl[2026], bl[2027], bl[2028], bl[2029], bl[2030], bl[2031], bl[2032], bl[2033], bl[2034], bl[2035], bl[2036], bl[2037], bl[2038], bl[2039], bl[2040], bl[2041], bl[2042], bl[2043], bl[2044], bl[2045], bl[2046], bl[2047], bl[2048], bl[2049], bl[2050], bl[2051], bl[2052], bl[2053], bl[2054], bl[2055], bl[2056], bl[2057], bl[2058], bl[2059], bl[2060], bl[2061], bl[2062], bl[2063], bl[2064], bl[2065], bl[2066], bl[2067], bl[2068], bl[2069], bl[2070], bl[2071], bl[2072], bl[2073], bl[2074], bl[2075], bl[2076], bl[2077], bl[2078], bl[2079], bl[2080], bl[2081], bl[2082], bl[2083], bl[2084], bl[2085], bl[2086], bl[2087], bl[2088], bl[2089], bl[2090], bl[2091], bl[2092], bl[2093], bl[2094], bl[2095], bl[2096], bl[2097], bl[2098], bl[2099], bl[2100], bl[2101], bl[2102], bl[2103], bl[2104], bl[2105], bl[2106], bl[2107], bl[2108], bl[2109], bl[2110], bl[2111], bl[2112], bl[2113], bl[2114], bl[2115], bl[2116], bl[2117], bl[2118], bl[2119], bl[2120], bl[2121], bl[2122], bl[2123], bl[2124], bl[2125], bl[2126], bl[2127], bl[2128], bl[2129], bl[2130], bl[2131], bl[2132], bl[2133], bl[2134], bl[2135], bl[2136], bl[2137], bl[2138], bl[2139], bl[2140], bl[2141], bl[2142], bl[2143], bl[2144], bl[2145], bl[2146], bl[2147], bl[2148], bl[2149], bl[2150], bl[2151], bl[2152], bl[2153], bl[2154], bl[2155], bl[2156], bl[2157], bl[2158], bl[2159], bl[2160], bl[2161], bl[2162], bl[2163], bl[2164], bl[2165], bl[2166], bl[2167], bl[2168], bl[2169], bl[2170], bl[2171], bl[2172], bl[2173], bl[2174], bl[2175], bl[2176], bl[2177], bl[2178], bl[2179], bl[2180], bl[2181], bl[2182], bl[2183], bl[2184], bl[2185], bl[2186], bl[2187], bl[2188], bl[2189], bl[2190], bl[2191], bl[2192], bl[2193], bl[2194], bl[2195], bl[2196], bl[2197], bl[2198], bl[2199], bl[2200], bl[2201], bl[2202], bl[2203], bl[2204], bl[2205], bl[2206], bl[2207], bl[2208], bl[2209], bl[2210], bl[2211], bl[2212], bl[2213], bl[2214], bl[2215], bl[2216], bl[2217], bl[2218], bl[2219], bl[2220], bl[2221], bl[2222], bl[2223], bl[2224], bl[2225], bl[2226], bl[2227], bl[2228], bl[2229], bl[2230], bl[2231], bl[2232], bl[2233], bl[2234], bl[2235], bl[2236], bl[2237], bl[2238], bl[2239], bl[2240], bl[2241], bl[2242], bl[2243], bl[2244], bl[2245], bl[2246], bl[2247], bl[2248], bl[2249], bl[2250], bl[2251], bl[2252], bl[2253], bl[2254], bl[2255], bl[2256], bl[2257], bl[2258], bl[2259], bl[2260], bl[2261], bl[2262], bl[2263], bl[2264], bl[2265], bl[2266], bl[2267], bl[2268], bl[2269], bl[2270], bl[2271], bl[2272], bl[2273], bl[2274], bl[2275], bl[2276], bl[2277], bl[2278], bl[2279], bl[2280], bl[2281], bl[2282], bl[2283], bl[2284], bl[2285], bl[2286], bl[2287], bl[2288], bl[2289], bl[2290], bl[2291], bl[2292], bl[2293], bl[2294], bl[2295], bl[2296], bl[2297], bl[2298], bl[2299], bl[2300], bl[2301], bl[2302], bl[2303], bl[2304], bl[2305], bl[2306], bl[2307], bl[2308], bl[2309], bl[2310], bl[2311], bl[2312], bl[2313], bl[2314], bl[2315], bl[2316], bl[2317], bl[2318], bl[2319], bl[2320], bl[2321], bl[2322], bl[2323], bl[2324], bl[2325], bl[2326], bl[2327], bl[2328], bl[2329], bl[2330], bl[2331], bl[2332], bl[2333], bl[2334], bl[2335], bl[2336], bl[2337], bl[2338], bl[2339], bl[2340], bl[2341], bl[2342], bl[2343], bl[2344], bl[2345], bl[2346], bl[2347], bl[2348], bl[2349], bl[2350], bl[2351], bl[2352], bl[2353], bl[2354], bl[2355], bl[2356], bl[2357], bl[2358], bl[2359], bl[2360], bl[2361], bl[2362], bl[2363], bl[2364], bl[2365], bl[2366], bl[2367], bl[2368], bl[2369], bl[2370], bl[2371], bl[2372], bl[2373], bl[2374], bl[2375], bl[2376], bl[2377], bl[2378], bl[2379], bl[2380], bl[2381], bl[2382], bl[2383], bl[2384], bl[2385], bl[2386], bl[2387], bl[2388], bl[2389], bl[2390], bl[2391], bl[2392], bl[2393], bl[2394], bl[2395], bl[2396], bl[2397], bl[2398], bl[2399], bl[2400], bl[2401], bl[2402], bl[2403], bl[2404], bl[2405], bl[2406], bl[2407], bl[2408], bl[2409], bl[2410], bl[2411], bl[2412], bl[2413], bl[2414], bl[2415], bl[2416], bl[2417], bl[2418], bl[2419], bl[2420], bl[2421], bl[2422], bl[2423], bl[2424], bl[2425], bl[2426], bl[2427], bl[2428], bl[2429], bl[2430], bl[2431], bl[2432], bl[2433], bl[2434], bl[2435], bl[2436], bl[2437], bl[2438], bl[2439], bl[2440], bl[2441], bl[2442], bl[2443], bl[2444], bl[2445], bl[2446], bl[2447], bl[2448], bl[2449], bl[2450], bl[2451], bl[2452], bl[2453], bl[2454], bl[2455], bl[2456], bl[2457], bl[2458], bl[2459], bl[2460], bl[2461], bl[2462], bl[2463], bl[2464], bl[2465], bl[2466], bl[2467], bl[2468], bl[2469], bl[2470], bl[2471], bl[2472], bl[2473], bl[2474], bl[2475], bl[2476], bl[2477], bl[2478], bl[2479], bl[2480], bl[2481], bl[2482], bl[2483], bl[2484], bl[2485], bl[2486], bl[2487], bl[2488], bl[2489], bl[2490], bl[2491], bl[2492], bl[2493], bl[2494], bl[2495], bl[2496], bl[2497], bl[2498], bl[2499], bl[2500], bl[2501], bl[2502], bl[2503], bl[2504], bl[2505], bl[2506], bl[2507], bl[2508], bl[2509], bl[2510], bl[2511], bl[2512], bl[2513], bl[2514], bl[2515], bl[2516], bl[2517], bl[2518], bl[2519], bl[2520], bl[2521], bl[2522], bl[2523], bl[2524], bl[2525], bl[2526], bl[2527], bl[2528], bl[2529], bl[2530], bl[2531], bl[2532], bl[2533], bl[2534], bl[2535], bl[2536], bl[2537], bl[2538], bl[2539], bl[2540], bl[2541], bl[2542], bl[2543], bl[2544], bl[2545], bl[2546], bl[2547], bl[2548], bl[2549], bl[2550], bl[2551], bl[2552], bl[2553], bl[2554], bl[2555], bl[2556], bl[2557], bl[2558], bl[2559], bl[2560], bl[2561], bl[2562], bl[2563], bl[2564], bl[2565], bl[2566], bl[2567], bl[2568], bl[2569], bl[2570], bl[2571], bl[2572], bl[2573], bl[2574], bl[2575], bl[2576], bl[2577], bl[2578], bl[2579], bl[2580], bl[2581], bl[2582], bl[2583], bl[2584], bl[2585], bl[2586], bl[2587], bl[2588], bl[2589], bl[2590], bl[2591], bl[2592], bl[2593], bl[2594], bl[2595], bl[2596], bl[2597], bl[2598], bl[2599], bl[2600], bl[2601], bl[2602], bl[2603], bl[2604], bl[2605], bl[2606], bl[2607], bl[2608], bl[2609], bl[2610], bl[2611], bl[2612], bl[2613], bl[2614], bl[2615], bl[2616], bl[2617], bl[2618], bl[2619], bl[2620], bl[2621], bl[2622], bl[2623], bl[2624], bl[2625], bl[2626], bl[2627], bl[2628], bl[2629], bl[2630], bl[2631], bl[2632], bl[2633], bl[2634], bl[2635], bl[2636], bl[2637], bl[2638], bl[2639], bl[2640], bl[2641], bl[2642], bl[2643], bl[2644], bl[2645], bl[2646], bl[2647], bl[2648], bl[2649], bl[2650], bl[2651], bl[2652], bl[2653], bl[2654], bl[2655], bl[2656], bl[2657], bl[2658], bl[2659], bl[2660], bl[2661], bl[2662], bl[2663], bl[2664], bl[2665], bl[2666], bl[2667], bl[10264], bl[10265], bl[10266], bl[10267], bl[10268], bl[10269], bl[10270], bl[10271], bl[10272], bl[10273], bl[10274], bl[10275], bl[10276], bl[10277], bl[10278], bl[10279], bl[10280], bl[10281], bl[10282], bl[10283], bl[10284], bl[10285], bl[10286], bl[10287], bl[10288], bl[10289], bl[10290], bl[10291], bl[10292], bl[10293], bl[10294], bl[10295], bl[10296], bl[10297], bl[10298], bl[10299], bl[10300], bl[10301], bl[10302], bl[10303], bl[10304], bl[10305], bl[10306], bl[10307], bl[10308], bl[10309], bl[10310], bl[10311], bl[10312], bl[10313], bl[10314], bl[10315], bl[10316], bl[10317], bl[10318], bl[10319], bl[10320], bl[10321], bl[10322], bl[10323], bl[10324], bl[10325], bl[10326], bl[10327], bl[10328], bl[10329], bl[10330], bl[10331], bl[10332], bl[10333], bl[10334], bl[10335], bl[10336], bl[10337], bl[10338], bl[10339], bl[10340], bl[10341], bl[10342], bl[10343], bl[1568], bl[1569], bl[1570], bl[1571], bl[1572], bl[1573], bl[1574], bl[1575], bl[1576], bl[1577], bl[1578], bl[1579], bl[1580], bl[1581], bl[1582], bl[1583], bl[1584], bl[1585], bl[1586], bl[1587], bl[1588], bl[1589], bl[1590], bl[1591], bl[1592], bl[1593], bl[1594], bl[1595], bl[1596], bl[1597], bl[1598], bl[1599], bl[1600], bl[1601], bl[1602], bl[1603], bl[1604], bl[1605], bl[1606], bl[1607], bl[1608], bl[1609], bl[1610], bl[1611], bl[1612], bl[1613], bl[1614], bl[1615], bl[1616], bl[1617], bl[1618], bl[1619], bl[1620], bl[1621], bl[1622], bl[1623], bl[1624], bl[1625], bl[1626], bl[1627], bl[1628], bl[1629], bl[1630], bl[1631], bl[1632], bl[1633], bl[1634], bl[1635], bl[1636], bl[1637], bl[1638], bl[1639], bl[1640], bl[1641], bl[1642], bl[1643], bl[1644], bl[1645], bl[1646], bl[1647], bl[10184], bl[10185], bl[10186], bl[10187], bl[10188], bl[10189], bl[10190], bl[10191], bl[10192], bl[10193], bl[10194], bl[10195], bl[10196], bl[10197], bl[10198], bl[10199], bl[10200], bl[10201], bl[10202], bl[10203], bl[10204], bl[10205], bl[10206], bl[10207], bl[10208], bl[10209], bl[10210], bl[10211], bl[10212], bl[10213], bl[10214], bl[10215], bl[10216], bl[10217], bl[10218], bl[10219], bl[10220], bl[10221], bl[10222], bl[10223], bl[10224], bl[10225], bl[10226], bl[10227], bl[10228], bl[10229], bl[10230], bl[10231], bl[10232], bl[10233], bl[10234], bl[10235], bl[10236], bl[10237], bl[10238], bl[10239], bl[10240], bl[10241], bl[10242], bl[10243], bl[10244], bl[10245], bl[10246], bl[10247], bl[10248], bl[10249], bl[10250], bl[10251], bl[10252], bl[10253], bl[10254], bl[10255], bl[10256], bl[10257], bl[10258], bl[10259], bl[10260], bl[10261], bl[10262], bl[10263]}),
        .wl({wl[1648], wl[1649], wl[1650], wl[1651], wl[1652], wl[1653], wl[1654], wl[1655], wl[1656], wl[1657], wl[1658], wl[1659], wl[1660], wl[1661], wl[1662], wl[1663], wl[1664], wl[1665], wl[1666], wl[1667], wl[1668], wl[1669], wl[1670], wl[1671], wl[1672], wl[1673], wl[1674], wl[1675], wl[1676], wl[1677], wl[1678], wl[1679], wl[1680], wl[1681], wl[1682], wl[1683], wl[1684], wl[1685], wl[1686], wl[1687], wl[1688], wl[1689], wl[1690], wl[1691], wl[1692], wl[1693], wl[1694], wl[1695], wl[1696], wl[1697], wl[1698], wl[1699], wl[1700], wl[1701], wl[1702], wl[1703], wl[1704], wl[1705], wl[1706], wl[1707], wl[1708], wl[1709], wl[1710], wl[1711], wl[1712], wl[1713], wl[1714], wl[1715], wl[1716], wl[1717], wl[1718], wl[1719], wl[1720], wl[1721], wl[1722], wl[1723], wl[1724], wl[1725], wl[1726], wl[1727], wl[1728], wl[1729], wl[1730], wl[1731], wl[1732], wl[1733], wl[1734], wl[1735], wl[1736], wl[1737], wl[1738], wl[1739], wl[1740], wl[1741], wl[1742], wl[1743], wl[1744], wl[1745], wl[1746], wl[1747], wl[1748], wl[1749], wl[1750], wl[1751], wl[1752], wl[1753], wl[1754], wl[1755], wl[1756], wl[1757], wl[1758], wl[1759], wl[1760], wl[1761], wl[1762], wl[1763], wl[1764], wl[1765], wl[1766], wl[1767], wl[1768], wl[1769], wl[1770], wl[1771], wl[1772], wl[1773], wl[1774], wl[1775], wl[1776], wl[1777], wl[1778], wl[1779], wl[1780], wl[1781], wl[1782], wl[1783], wl[1784], wl[1785], wl[1786], wl[1787], wl[1788], wl[1789], wl[1790], wl[1791], wl[1792], wl[1793], wl[1794], wl[1795], wl[1796], wl[1797], wl[1798], wl[1799], wl[1800], wl[1801], wl[1802], wl[1803], wl[1804], wl[1805], wl[1806], wl[1807], wl[1808], wl[1809], wl[1810], wl[1811], wl[1812], wl[1813], wl[1814], wl[1815], wl[1816], wl[1817], wl[1818], wl[1819], wl[1820], wl[1821], wl[1822], wl[1823], wl[1824], wl[1825], wl[1826], wl[1827], wl[1828], wl[1829], wl[1830], wl[1831], wl[1832], wl[1833], wl[1834], wl[1835], wl[1836], wl[1837], wl[1838], wl[1839], wl[1840], wl[1841], wl[1842], wl[1843], wl[1844], wl[1845], wl[1846], wl[1847], wl[1848], wl[1849], wl[1850], wl[1851], wl[1852], wl[1853], wl[1854], wl[1855], wl[1856], wl[1857], wl[1858], wl[1859], wl[1860], wl[1861], wl[1862], wl[1863], wl[1864], wl[1865], wl[1866], wl[1867], wl[1868], wl[1869], wl[1870], wl[1871], wl[1872], wl[1873], wl[1874], wl[1875], wl[1876], wl[1877], wl[1878], wl[1879], wl[1880], wl[1881], wl[1882], wl[1883], wl[1884], wl[1885], wl[1886], wl[1887], wl[1888], wl[1889], wl[1890], wl[1891], wl[1892], wl[1893], wl[1894], wl[1895], wl[1896], wl[1897], wl[1898], wl[1899], wl[1900], wl[1901], wl[1902], wl[1903], wl[1904], wl[1905], wl[1906], wl[1907], wl[1908], wl[1909], wl[1910], wl[1911], wl[1912], wl[1913], wl[1914], wl[1915], wl[1916], wl[1917], wl[1918], wl[1919], wl[1920], wl[1921], wl[1922], wl[1923], wl[1924], wl[1925], wl[1926], wl[1927], wl[1928], wl[1929], wl[1930], wl[1931], wl[1932], wl[1933], wl[1934], wl[1935], wl[1936], wl[1937], wl[1938], wl[1939], wl[1940], wl[1941], wl[1942], wl[1943], wl[1944], wl[1945], wl[1946], wl[1947], wl[1948], wl[1949], wl[1950], wl[1951], wl[1952], wl[1953], wl[1954], wl[1955], wl[1956], wl[1957], wl[1958], wl[1959], wl[1960], wl[1961], wl[1962], wl[1963], wl[1964], wl[1965], wl[1966], wl[1967], wl[1968], wl[1969], wl[1970], wl[1971], wl[1972], wl[1973], wl[1974], wl[1975], wl[1976], wl[1977], wl[1978], wl[1979], wl[1980], wl[1981], wl[1982], wl[1983], wl[1984], wl[1985], wl[1986], wl[1987], wl[1988], wl[1989], wl[1990], wl[1991], wl[1992], wl[1993], wl[1994], wl[1995], wl[1996], wl[1997], wl[1998], wl[1999], wl[2000], wl[2001], wl[2002], wl[2003], wl[2004], wl[2005], wl[2006], wl[2007], wl[2008], wl[2009], wl[2010], wl[2011], wl[2012], wl[2013], wl[2014], wl[2015], wl[2016], wl[2017], wl[2018], wl[2019], wl[2020], wl[2021], wl[2022], wl[2023], wl[2024], wl[2025], wl[2026], wl[2027], wl[2028], wl[2029], wl[2030], wl[2031], wl[2032], wl[2033], wl[2034], wl[2035], wl[2036], wl[2037], wl[2038], wl[2039], wl[2040], wl[2041], wl[2042], wl[2043], wl[2044], wl[2045], wl[2046], wl[2047], wl[2048], wl[2049], wl[2050], wl[2051], wl[2052], wl[2053], wl[2054], wl[2055], wl[2056], wl[2057], wl[2058], wl[2059], wl[2060], wl[2061], wl[2062], wl[2063], wl[2064], wl[2065], wl[2066], wl[2067], wl[2068], wl[2069], wl[2070], wl[2071], wl[2072], wl[2073], wl[2074], wl[2075], wl[2076], wl[2077], wl[2078], wl[2079], wl[2080], wl[2081], wl[2082], wl[2083], wl[2084], wl[2085], wl[2086], wl[2087], wl[2088], wl[2089], wl[2090], wl[2091], wl[2092], wl[2093], wl[2094], wl[2095], wl[2096], wl[2097], wl[2098], wl[2099], wl[2100], wl[2101], wl[2102], wl[2103], wl[2104], wl[2105], wl[2106], wl[2107], wl[2108], wl[2109], wl[2110], wl[2111], wl[2112], wl[2113], wl[2114], wl[2115], wl[2116], wl[2117], wl[2118], wl[2119], wl[2120], wl[2121], wl[2122], wl[2123], wl[2124], wl[2125], wl[2126], wl[2127], wl[2128], wl[2129], wl[2130], wl[2131], wl[2132], wl[2133], wl[2134], wl[2135], wl[2136], wl[2137], wl[2138], wl[2139], wl[2140], wl[2141], wl[2142], wl[2143], wl[2144], wl[2145], wl[2146], wl[2147], wl[2148], wl[2149], wl[2150], wl[2151], wl[2152], wl[2153], wl[2154], wl[2155], wl[2156], wl[2157], wl[2158], wl[2159], wl[2160], wl[2161], wl[2162], wl[2163], wl[2164], wl[2165], wl[2166], wl[2167], wl[2168], wl[2169], wl[2170], wl[2171], wl[2172], wl[2173], wl[2174], wl[2175], wl[2176], wl[2177], wl[2178], wl[2179], wl[2180], wl[2181], wl[2182], wl[2183], wl[2184], wl[2185], wl[2186], wl[2187], wl[2188], wl[2189], wl[2190], wl[2191], wl[2192], wl[2193], wl[2194], wl[2195], wl[2196], wl[2197], wl[2198], wl[2199], wl[2200], wl[2201], wl[2202], wl[2203], wl[2204], wl[2205], wl[2206], wl[2207], wl[2208], wl[2209], wl[2210], wl[2211], wl[2212], wl[2213], wl[2214], wl[2215], wl[2216], wl[2217], wl[2218], wl[2219], wl[2220], wl[2221], wl[2222], wl[2223], wl[2224], wl[2225], wl[2226], wl[2227], wl[2228], wl[2229], wl[2230], wl[2231], wl[2232], wl[2233], wl[2234], wl[2235], wl[2236], wl[2237], wl[2238], wl[2239], wl[2240], wl[2241], wl[2242], wl[2243], wl[2244], wl[2245], wl[2246], wl[2247], wl[2248], wl[2249], wl[2250], wl[2251], wl[2252], wl[2253], wl[2254], wl[2255], wl[2256], wl[2257], wl[2258], wl[2259], wl[2260], wl[2261], wl[2262], wl[2263], wl[2264], wl[2265], wl[2266], wl[2267], wl[2268], wl[2269], wl[2270], wl[2271], wl[2272], wl[2273], wl[2274], wl[2275], wl[2276], wl[2277], wl[2278], wl[2279], wl[2280], wl[2281], wl[2282], wl[2283], wl[2284], wl[2285], wl[2286], wl[2287], wl[2288], wl[2289], wl[2290], wl[2291], wl[2292], wl[2293], wl[2294], wl[2295], wl[2296], wl[2297], wl[2298], wl[2299], wl[2300], wl[2301], wl[2302], wl[2303], wl[2304], wl[2305], wl[2306], wl[2307], wl[2308], wl[2309], wl[2310], wl[2311], wl[2312], wl[2313], wl[2314], wl[2315], wl[2316], wl[2317], wl[2318], wl[2319], wl[2320], wl[2321], wl[2322], wl[2323], wl[2324], wl[2325], wl[2326], wl[2327], wl[2328], wl[2329], wl[2330], wl[2331], wl[2332], wl[2333], wl[2334], wl[2335], wl[2336], wl[2337], wl[2338], wl[2339], wl[2340], wl[2341], wl[2342], wl[2343], wl[2344], wl[2345], wl[2346], wl[2347], wl[2348], wl[2349], wl[2350], wl[2351], wl[2352], wl[2353], wl[2354], wl[2355], wl[2356], wl[2357], wl[2358], wl[2359], wl[2360], wl[2361], wl[2362], wl[2363], wl[2364], wl[2365], wl[2366], wl[2367], wl[2368], wl[2369], wl[2370], wl[2371], wl[2372], wl[2373], wl[2374], wl[2375], wl[2376], wl[2377], wl[2378], wl[2379], wl[2380], wl[2381], wl[2382], wl[2383], wl[2384], wl[2385], wl[2386], wl[2387], wl[2388], wl[2389], wl[2390], wl[2391], wl[2392], wl[2393], wl[2394], wl[2395], wl[2396], wl[2397], wl[2398], wl[2399], wl[2400], wl[2401], wl[2402], wl[2403], wl[2404], wl[2405], wl[2406], wl[2407], wl[2408], wl[2409], wl[2410], wl[2411], wl[2412], wl[2413], wl[2414], wl[2415], wl[2416], wl[2417], wl[2418], wl[2419], wl[2420], wl[2421], wl[2422], wl[2423], wl[2424], wl[2425], wl[2426], wl[2427], wl[2428], wl[2429], wl[2430], wl[2431], wl[2432], wl[2433], wl[2434], wl[2435], wl[2436], wl[2437], wl[2438], wl[2439], wl[2440], wl[2441], wl[2442], wl[2443], wl[2444], wl[2445], wl[2446], wl[2447], wl[2448], wl[2449], wl[2450], wl[2451], wl[2452], wl[2453], wl[2454], wl[2455], wl[2456], wl[2457], wl[2458], wl[2459], wl[2460], wl[2461], wl[2462], wl[2463], wl[2464], wl[2465], wl[2466], wl[2467], wl[2468], wl[2469], wl[2470], wl[2471], wl[2472], wl[2473], wl[2474], wl[2475], wl[2476], wl[2477], wl[2478], wl[2479], wl[2480], wl[2481], wl[2482], wl[2483], wl[2484], wl[2485], wl[2486], wl[2487], wl[2488], wl[2489], wl[2490], wl[2491], wl[2492], wl[2493], wl[2494], wl[2495], wl[2496], wl[2497], wl[2498], wl[2499], wl[2500], wl[2501], wl[2502], wl[2503], wl[2504], wl[2505], wl[2506], wl[2507], wl[2508], wl[2509], wl[2510], wl[2511], wl[2512], wl[2513], wl[2514], wl[2515], wl[2516], wl[2517], wl[2518], wl[2519], wl[2520], wl[2521], wl[2522], wl[2523], wl[2524], wl[2525], wl[2526], wl[2527], wl[2528], wl[2529], wl[2530], wl[2531], wl[2532], wl[2533], wl[2534], wl[2535], wl[2536], wl[2537], wl[2538], wl[2539], wl[2540], wl[2541], wl[2542], wl[2543], wl[2544], wl[2545], wl[2546], wl[2547], wl[2548], wl[2549], wl[2550], wl[2551], wl[2552], wl[2553], wl[2554], wl[2555], wl[2556], wl[2557], wl[2558], wl[2559], wl[2560], wl[2561], wl[2562], wl[2563], wl[2564], wl[2565], wl[2566], wl[2567], wl[2568], wl[2569], wl[2570], wl[2571], wl[2572], wl[2573], wl[2574], wl[2575], wl[2576], wl[2577], wl[2578], wl[2579], wl[2580], wl[2581], wl[2582], wl[2583], wl[2584], wl[2585], wl[2586], wl[2587], wl[2588], wl[2589], wl[2590], wl[2591], wl[2592], wl[2593], wl[2594], wl[2595], wl[2596], wl[2597], wl[2598], wl[2599], wl[2600], wl[2601], wl[2602], wl[2603], wl[2604], wl[2605], wl[2606], wl[2607], wl[2608], wl[2609], wl[2610], wl[2611], wl[2612], wl[2613], wl[2614], wl[2615], wl[2616], wl[2617], wl[2618], wl[2619], wl[2620], wl[2621], wl[2622], wl[2623], wl[2624], wl[2625], wl[2626], wl[2627], wl[2628], wl[2629], wl[2630], wl[2631], wl[2632], wl[2633], wl[2634], wl[2635], wl[2636], wl[2637], wl[2638], wl[2639], wl[2640], wl[2641], wl[2642], wl[2643], wl[2644], wl[2645], wl[2646], wl[2647], wl[2648], wl[2649], wl[2650], wl[2651], wl[2652], wl[2653], wl[2654], wl[2655], wl[2656], wl[2657], wl[2658], wl[2659], wl[2660], wl[2661], wl[2662], wl[2663], wl[2664], wl[2665], wl[2666], wl[2667], wl[10264], wl[10265], wl[10266], wl[10267], wl[10268], wl[10269], wl[10270], wl[10271], wl[10272], wl[10273], wl[10274], wl[10275], wl[10276], wl[10277], wl[10278], wl[10279], wl[10280], wl[10281], wl[10282], wl[10283], wl[10284], wl[10285], wl[10286], wl[10287], wl[10288], wl[10289], wl[10290], wl[10291], wl[10292], wl[10293], wl[10294], wl[10295], wl[10296], wl[10297], wl[10298], wl[10299], wl[10300], wl[10301], wl[10302], wl[10303], wl[10304], wl[10305], wl[10306], wl[10307], wl[10308], wl[10309], wl[10310], wl[10311], wl[10312], wl[10313], wl[10314], wl[10315], wl[10316], wl[10317], wl[10318], wl[10319], wl[10320], wl[10321], wl[10322], wl[10323], wl[10324], wl[10325], wl[10326], wl[10327], wl[10328], wl[10329], wl[10330], wl[10331], wl[10332], wl[10333], wl[10334], wl[10335], wl[10336], wl[10337], wl[10338], wl[10339], wl[10340], wl[10341], wl[10342], wl[10343], wl[1568], wl[1569], wl[1570], wl[1571], wl[1572], wl[1573], wl[1574], wl[1575], wl[1576], wl[1577], wl[1578], wl[1579], wl[1580], wl[1581], wl[1582], wl[1583], wl[1584], wl[1585], wl[1586], wl[1587], wl[1588], wl[1589], wl[1590], wl[1591], wl[1592], wl[1593], wl[1594], wl[1595], wl[1596], wl[1597], wl[1598], wl[1599], wl[1600], wl[1601], wl[1602], wl[1603], wl[1604], wl[1605], wl[1606], wl[1607], wl[1608], wl[1609], wl[1610], wl[1611], wl[1612], wl[1613], wl[1614], wl[1615], wl[1616], wl[1617], wl[1618], wl[1619], wl[1620], wl[1621], wl[1622], wl[1623], wl[1624], wl[1625], wl[1626], wl[1627], wl[1628], wl[1629], wl[1630], wl[1631], wl[1632], wl[1633], wl[1634], wl[1635], wl[1636], wl[1637], wl[1638], wl[1639], wl[1640], wl[1641], wl[1642], wl[1643], wl[1644], wl[1645], wl[1646], wl[1647], wl[10184], wl[10185], wl[10186], wl[10187], wl[10188], wl[10189], wl[10190], wl[10191], wl[10192], wl[10193], wl[10194], wl[10195], wl[10196], wl[10197], wl[10198], wl[10199], wl[10200], wl[10201], wl[10202], wl[10203], wl[10204], wl[10205], wl[10206], wl[10207], wl[10208], wl[10209], wl[10210], wl[10211], wl[10212], wl[10213], wl[10214], wl[10215], wl[10216], wl[10217], wl[10218], wl[10219], wl[10220], wl[10221], wl[10222], wl[10223], wl[10224], wl[10225], wl[10226], wl[10227], wl[10228], wl[10229], wl[10230], wl[10231], wl[10232], wl[10233], wl[10234], wl[10235], wl[10236], wl[10237], wl[10238], wl[10239], wl[10240], wl[10241], wl[10242], wl[10243], wl[10244], wl[10245], wl[10246], wl[10247], wl[10248], wl[10249], wl[10250], wl[10251], wl[10252], wl[10253], wl[10254], wl[10255], wl[10256], wl[10257], wl[10258], wl[10259], wl[10260], wl[10261], wl[10262], wl[10263]})
    );
    tile tile_2__3_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_0__2__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_0__2__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_0__2__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_1__1__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_1__1__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_1__1__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_0__1__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_0__1__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_0__1__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_0__1__grid_top_r_in[1]),
        .grid_left_in(grid_clb_1__2__grid_left_in),
        .grid_bottom_in(grid_clb_1__2__grid_bottom_in),
        .chanx_left_in(sb_0__1__1_chanx_right_out),
        .chanx_left_out(cbx_1__1__1_chanx_left_out),
        .grid_top_out(grid_clb_1__3__grid_bottom_in),
        .chany_bottom_in(sb_1__1__0_chany_top_out),
        .chany_bottom_out(cby_1__1__1_chany_bottom_out),
        .grid_right_out(grid_clb_2__2__grid_left_in),
        .chany_top_in_0(cby_1__1__2_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__4_chanx_left_out),
        .chany_top_out_0(sb_1__1__1_chany_top_out),
        .chanx_right_out_0(sb_1__1__1_chanx_right_out),
        .grid_top_r_in(sb_1__2__grid_top_r_in),
        .grid_top_l_in(sb_1__2__grid_top_l_in),
        .grid_right_t_in(sb_1__2__grid_right_t_in),
        .grid_right_b_in(sb_1__2__grid_right_b_in),
        .grid_bottom_r_in(sb_1__1__grid_top_r_in),
        .grid_bottom_l_in(sb_1__1__grid_top_l_in),
        .grid_left_t_in(sb_0__2__grid_right_t_in),
        .grid_left_b_in(sb_0__2__grid_right_b_in),
        .bl({bl[10424], bl[10425], bl[10426], bl[10427], bl[10428], bl[10429], bl[10430], bl[10431], bl[10432], bl[10433], bl[10434], bl[10435], bl[10436], bl[10437], bl[10438], bl[10439], bl[10440], bl[10441], bl[10442], bl[10443], bl[10444], bl[10445], bl[10446], bl[10447], bl[10448], bl[10449], bl[10450], bl[10451], bl[10452], bl[10453], bl[10454], bl[10455], bl[10456], bl[10457], bl[10458], bl[10459], bl[10460], bl[10461], bl[10462], bl[10463], bl[10464], bl[10465], bl[10466], bl[10467], bl[10468], bl[10469], bl[10470], bl[10471], bl[10472], bl[10473], bl[10474], bl[10475], bl[10476], bl[10477], bl[10478], bl[10479], bl[10480], bl[10481], bl[10482], bl[10483], bl[10484], bl[10485], bl[10486], bl[10487], bl[10488], bl[10489], bl[10490], bl[10491], bl[10492], bl[10493], bl[10494], bl[10495], bl[10496], bl[10497], bl[10498], bl[10499], bl[10500], bl[10501], bl[10502], bl[10503], bl[10504], bl[10505], bl[10506], bl[10507], bl[10508], bl[10509], bl[10510], bl[10511], bl[10512], bl[10513], bl[10514], bl[10515], bl[10516], bl[10517], bl[10518], bl[10519], bl[10520], bl[10521], bl[10522], bl[10523], bl[10524], bl[10525], bl[10526], bl[10527], bl[10528], bl[10529], bl[10530], bl[10531], bl[10532], bl[10533], bl[10534], bl[10535], bl[10536], bl[10537], bl[10538], bl[10539], bl[10540], bl[10541], bl[10542], bl[10543], bl[10544], bl[10545], bl[10546], bl[10547], bl[10548], bl[10549], bl[10550], bl[10551], bl[10552], bl[10553], bl[10554], bl[10555], bl[10556], bl[10557], bl[10558], bl[10559], bl[10560], bl[10561], bl[10562], bl[10563], bl[10564], bl[10565], bl[10566], bl[10567], bl[10568], bl[10569], bl[10570], bl[10571], bl[10572], bl[10573], bl[10574], bl[10575], bl[10576], bl[10577], bl[10578], bl[10579], bl[10580], bl[10581], bl[10582], bl[10583], bl[10584], bl[10585], bl[10586], bl[10587], bl[10588], bl[10589], bl[10590], bl[10591], bl[10592], bl[10593], bl[10594], bl[10595], bl[10596], bl[10597], bl[10598], bl[10599], bl[10600], bl[10601], bl[10602], bl[10603], bl[10604], bl[10605], bl[10606], bl[10607], bl[10608], bl[10609], bl[10610], bl[10611], bl[10612], bl[10613], bl[10614], bl[10615], bl[10616], bl[10617], bl[10618], bl[10619], bl[10620], bl[10621], bl[10622], bl[10623], bl[10624], bl[10625], bl[10626], bl[10627], bl[10628], bl[10629], bl[10630], bl[10631], bl[10632], bl[10633], bl[10634], bl[10635], bl[10636], bl[10637], bl[10638], bl[10639], bl[10640], bl[10641], bl[10642], bl[10643], bl[10644], bl[10645], bl[10646], bl[10647], bl[10648], bl[10649], bl[10650], bl[10651], bl[10652], bl[10653], bl[10654], bl[10655], bl[10656], bl[10657], bl[10658], bl[10659], bl[10660], bl[10661], bl[10662], bl[10663], bl[10664], bl[10665], bl[10666], bl[10667], bl[10668], bl[10669], bl[10670], bl[10671], bl[10672], bl[10673], bl[10674], bl[10675], bl[10676], bl[10677], bl[10678], bl[10679], bl[10680], bl[10681], bl[10682], bl[10683], bl[10684], bl[10685], bl[10686], bl[10687], bl[10688], bl[10689], bl[10690], bl[10691], bl[10692], bl[10693], bl[10694], bl[10695], bl[10696], bl[10697], bl[10698], bl[10699], bl[10700], bl[10701], bl[10702], bl[10703], bl[10704], bl[10705], bl[10706], bl[10707], bl[10708], bl[10709], bl[10710], bl[10711], bl[10712], bl[10713], bl[10714], bl[10715], bl[10716], bl[10717], bl[10718], bl[10719], bl[10720], bl[10721], bl[10722], bl[10723], bl[10724], bl[10725], bl[10726], bl[10727], bl[10728], bl[10729], bl[10730], bl[10731], bl[10732], bl[10733], bl[10734], bl[10735], bl[10736], bl[10737], bl[10738], bl[10739], bl[10740], bl[10741], bl[10742], bl[10743], bl[10744], bl[10745], bl[10746], bl[10747], bl[10748], bl[10749], bl[10750], bl[10751], bl[10752], bl[10753], bl[10754], bl[10755], bl[10756], bl[10757], bl[10758], bl[10759], bl[10760], bl[10761], bl[10762], bl[10763], bl[10764], bl[10765], bl[10766], bl[10767], bl[10768], bl[10769], bl[10770], bl[10771], bl[10772], bl[10773], bl[10774], bl[10775], bl[10776], bl[10777], bl[10778], bl[10779], bl[10780], bl[10781], bl[10782], bl[10783], bl[10784], bl[10785], bl[10786], bl[10787], bl[10788], bl[10789], bl[10790], bl[10791], bl[10792], bl[10793], bl[10794], bl[10795], bl[10796], bl[10797], bl[10798], bl[10799], bl[10800], bl[10801], bl[10802], bl[10803], bl[10804], bl[10805], bl[10806], bl[10807], bl[10808], bl[10809], bl[10810], bl[10811], bl[10812], bl[10813], bl[10814], bl[10815], bl[10816], bl[10817], bl[10818], bl[10819], bl[10820], bl[10821], bl[10822], bl[10823], bl[10824], bl[10825], bl[10826], bl[10827], bl[10828], bl[10829], bl[10830], bl[10831], bl[10832], bl[10833], bl[10834], bl[10835], bl[10836], bl[10837], bl[10838], bl[10839], bl[10840], bl[10841], bl[10842], bl[10843], bl[10844], bl[10845], bl[10846], bl[10847], bl[10848], bl[10849], bl[10850], bl[10851], bl[10852], bl[10853], bl[10854], bl[10855], bl[10856], bl[10857], bl[10858], bl[10859], bl[10860], bl[10861], bl[10862], bl[10863], bl[10864], bl[10865], bl[10866], bl[10867], bl[10868], bl[10869], bl[10870], bl[10871], bl[10872], bl[10873], bl[10874], bl[10875], bl[10876], bl[10877], bl[10878], bl[10879], bl[10880], bl[10881], bl[10882], bl[10883], bl[10884], bl[10885], bl[10886], bl[10887], bl[10888], bl[10889], bl[10890], bl[10891], bl[10892], bl[10893], bl[10894], bl[10895], bl[10896], bl[10897], bl[10898], bl[10899], bl[10900], bl[10901], bl[10902], bl[10903], bl[10904], bl[10905], bl[10906], bl[10907], bl[10908], bl[10909], bl[10910], bl[10911], bl[10912], bl[10913], bl[10914], bl[10915], bl[10916], bl[10917], bl[10918], bl[10919], bl[10920], bl[10921], bl[10922], bl[10923], bl[10924], bl[10925], bl[10926], bl[10927], bl[10928], bl[10929], bl[10930], bl[10931], bl[10932], bl[10933], bl[10934], bl[10935], bl[10936], bl[10937], bl[10938], bl[10939], bl[10940], bl[10941], bl[10942], bl[10943], bl[10944], bl[10945], bl[10946], bl[10947], bl[10948], bl[10949], bl[10950], bl[10951], bl[10952], bl[10953], bl[10954], bl[10955], bl[10956], bl[10957], bl[10958], bl[10959], bl[10960], bl[10961], bl[10962], bl[10963], bl[10964], bl[10965], bl[10966], bl[10967], bl[10968], bl[10969], bl[10970], bl[10971], bl[10972], bl[10973], bl[10974], bl[10975], bl[10976], bl[10977], bl[10978], bl[10979], bl[10980], bl[10981], bl[10982], bl[10983], bl[10984], bl[10985], bl[10986], bl[10987], bl[10988], bl[10989], bl[10990], bl[10991], bl[10992], bl[10993], bl[10994], bl[10995], bl[10996], bl[10997], bl[10998], bl[10999], bl[11000], bl[11001], bl[11002], bl[11003], bl[11004], bl[11005], bl[11006], bl[11007], bl[11008], bl[11009], bl[11010], bl[11011], bl[11012], bl[11013], bl[11014], bl[11015], bl[11016], bl[11017], bl[11018], bl[11019], bl[11020], bl[11021], bl[11022], bl[11023], bl[11024], bl[11025], bl[11026], bl[11027], bl[11028], bl[11029], bl[11030], bl[11031], bl[11032], bl[11033], bl[11034], bl[11035], bl[11036], bl[11037], bl[11038], bl[11039], bl[11040], bl[11041], bl[11042], bl[11043], bl[11044], bl[11045], bl[11046], bl[11047], bl[11048], bl[11049], bl[11050], bl[11051], bl[11052], bl[11053], bl[11054], bl[11055], bl[11056], bl[11057], bl[11058], bl[11059], bl[11060], bl[11061], bl[11062], bl[11063], bl[11064], bl[11065], bl[11066], bl[11067], bl[11068], bl[11069], bl[11070], bl[11071], bl[11072], bl[11073], bl[11074], bl[11075], bl[11076], bl[11077], bl[11078], bl[11079], bl[11080], bl[11081], bl[11082], bl[11083], bl[11084], bl[11085], bl[11086], bl[11087], bl[11088], bl[11089], bl[11090], bl[11091], bl[11092], bl[11093], bl[11094], bl[11095], bl[11096], bl[11097], bl[11098], bl[11099], bl[11100], bl[11101], bl[11102], bl[11103], bl[11104], bl[11105], bl[11106], bl[11107], bl[11108], bl[11109], bl[11110], bl[11111], bl[11112], bl[11113], bl[11114], bl[11115], bl[11116], bl[11117], bl[11118], bl[11119], bl[11120], bl[11121], bl[11122], bl[11123], bl[11124], bl[11125], bl[11126], bl[11127], bl[11128], bl[11129], bl[11130], bl[11131], bl[11132], bl[11133], bl[11134], bl[11135], bl[11136], bl[11137], bl[11138], bl[11139], bl[11140], bl[11141], bl[11142], bl[11143], bl[11144], bl[11145], bl[11146], bl[11147], bl[11148], bl[11149], bl[11150], bl[11151], bl[11152], bl[11153], bl[11154], bl[11155], bl[11156], bl[11157], bl[11158], bl[11159], bl[11160], bl[11161], bl[11162], bl[11163], bl[11164], bl[11165], bl[11166], bl[11167], bl[11168], bl[11169], bl[11170], bl[11171], bl[11172], bl[11173], bl[11174], bl[11175], bl[11176], bl[11177], bl[11178], bl[11179], bl[11180], bl[11181], bl[11182], bl[11183], bl[11184], bl[11185], bl[11186], bl[11187], bl[11188], bl[11189], bl[11190], bl[11191], bl[11192], bl[11193], bl[11194], bl[11195], bl[11196], bl[11197], bl[11198], bl[11199], bl[11200], bl[11201], bl[11202], bl[11203], bl[11204], bl[11205], bl[11206], bl[11207], bl[11208], bl[11209], bl[11210], bl[11211], bl[11212], bl[11213], bl[11214], bl[11215], bl[11216], bl[11217], bl[11218], bl[11219], bl[11220], bl[11221], bl[11222], bl[11223], bl[11224], bl[11225], bl[11226], bl[11227], bl[11228], bl[11229], bl[11230], bl[11231], bl[11232], bl[11233], bl[11234], bl[11235], bl[11236], bl[11237], bl[11238], bl[11239], bl[11240], bl[11241], bl[11242], bl[11243], bl[11244], bl[11245], bl[11246], bl[11247], bl[11248], bl[11249], bl[11250], bl[11251], bl[11252], bl[11253], bl[11254], bl[11255], bl[11256], bl[11257], bl[11258], bl[11259], bl[11260], bl[11261], bl[11262], bl[11263], bl[11264], bl[11265], bl[11266], bl[11267], bl[11268], bl[11269], bl[11270], bl[11271], bl[11272], bl[11273], bl[11274], bl[11275], bl[11276], bl[11277], bl[11278], bl[11279], bl[11280], bl[11281], bl[11282], bl[11283], bl[11284], bl[11285], bl[11286], bl[11287], bl[11288], bl[11289], bl[11290], bl[11291], bl[11292], bl[11293], bl[11294], bl[11295], bl[11296], bl[11297], bl[11298], bl[11299], bl[11300], bl[11301], bl[11302], bl[11303], bl[11304], bl[11305], bl[11306], bl[11307], bl[11308], bl[11309], bl[11310], bl[11311], bl[11312], bl[11313], bl[11314], bl[11315], bl[11316], bl[11317], bl[11318], bl[11319], bl[11320], bl[11321], bl[11322], bl[11323], bl[11324], bl[11325], bl[11326], bl[11327], bl[11328], bl[11329], bl[11330], bl[11331], bl[11332], bl[11333], bl[11334], bl[11335], bl[11336], bl[11337], bl[11338], bl[11339], bl[11340], bl[11341], bl[11342], bl[11343], bl[11344], bl[11345], bl[11346], bl[11347], bl[11348], bl[11349], bl[11350], bl[11351], bl[11352], bl[11353], bl[11354], bl[11355], bl[11356], bl[11357], bl[11358], bl[11359], bl[11360], bl[11361], bl[11362], bl[11363], bl[11364], bl[11365], bl[11366], bl[11367], bl[11368], bl[11369], bl[11370], bl[11371], bl[11372], bl[11373], bl[11374], bl[11375], bl[11376], bl[11377], bl[11378], bl[11379], bl[11380], bl[11381], bl[11382], bl[11383], bl[11384], bl[11385], bl[11386], bl[11387], bl[11388], bl[11389], bl[11390], bl[11391], bl[11392], bl[11393], bl[11394], bl[11395], bl[11396], bl[11397], bl[11398], bl[11399], bl[11400], bl[11401], bl[11402], bl[11403], bl[11404], bl[11405], bl[11406], bl[11407], bl[11408], bl[11409], bl[11410], bl[11411], bl[11412], bl[11413], bl[11414], bl[11415], bl[11416], bl[11417], bl[11418], bl[11419], bl[11420], bl[11421], bl[11422], bl[11423], bl[11424], bl[11425], bl[11426], bl[11427], bl[11428], bl[11429], bl[11430], bl[11431], bl[11432], bl[11433], bl[11434], bl[11435], bl[11436], bl[11437], bl[11438], bl[11439], bl[11440], bl[11441], bl[11442], bl[11443], bl[11524], bl[11525], bl[11526], bl[11527], bl[11528], bl[11529], bl[11530], bl[11531], bl[11532], bl[11533], bl[11534], bl[11535], bl[11536], bl[11537], bl[11538], bl[11539], bl[11540], bl[11541], bl[11542], bl[11543], bl[11544], bl[11545], bl[11546], bl[11547], bl[11548], bl[11549], bl[11550], bl[11551], bl[11552], bl[11553], bl[11554], bl[11555], bl[11556], bl[11557], bl[11558], bl[11559], bl[11560], bl[11561], bl[11562], bl[11563], bl[11564], bl[11565], bl[11566], bl[11567], bl[11568], bl[11569], bl[11570], bl[11571], bl[11572], bl[11573], bl[11574], bl[11575], bl[11576], bl[11577], bl[11578], bl[11579], bl[11580], bl[11581], bl[11582], bl[11583], bl[11584], bl[11585], bl[11586], bl[11587], bl[11588], bl[11589], bl[11590], bl[11591], bl[11592], bl[11593], bl[11594], bl[11595], bl[11596], bl[11597], bl[11598], bl[11599], bl[11600], bl[11601], bl[11602], bl[11603], bl[10344], bl[10345], bl[10346], bl[10347], bl[10348], bl[10349], bl[10350], bl[10351], bl[10352], bl[10353], bl[10354], bl[10355], bl[10356], bl[10357], bl[10358], bl[10359], bl[10360], bl[10361], bl[10362], bl[10363], bl[10364], bl[10365], bl[10366], bl[10367], bl[10368], bl[10369], bl[10370], bl[10371], bl[10372], bl[10373], bl[10374], bl[10375], bl[10376], bl[10377], bl[10378], bl[10379], bl[10380], bl[10381], bl[10382], bl[10383], bl[10384], bl[10385], bl[10386], bl[10387], bl[10388], bl[10389], bl[10390], bl[10391], bl[10392], bl[10393], bl[10394], bl[10395], bl[10396], bl[10397], bl[10398], bl[10399], bl[10400], bl[10401], bl[10402], bl[10403], bl[10404], bl[10405], bl[10406], bl[10407], bl[10408], bl[10409], bl[10410], bl[10411], bl[10412], bl[10413], bl[10414], bl[10415], bl[10416], bl[10417], bl[10418], bl[10419], bl[10420], bl[10421], bl[10422], bl[10423], bl[11444], bl[11445], bl[11446], bl[11447], bl[11448], bl[11449], bl[11450], bl[11451], bl[11452], bl[11453], bl[11454], bl[11455], bl[11456], bl[11457], bl[11458], bl[11459], bl[11460], bl[11461], bl[11462], bl[11463], bl[11464], bl[11465], bl[11466], bl[11467], bl[11468], bl[11469], bl[11470], bl[11471], bl[11472], bl[11473], bl[11474], bl[11475], bl[11476], bl[11477], bl[11478], bl[11479], bl[11480], bl[11481], bl[11482], bl[11483], bl[11484], bl[11485], bl[11486], bl[11487], bl[11488], bl[11489], bl[11490], bl[11491], bl[11492], bl[11493], bl[11494], bl[11495], bl[11496], bl[11497], bl[11498], bl[11499], bl[11500], bl[11501], bl[11502], bl[11503], bl[11504], bl[11505], bl[11506], bl[11507], bl[11508], bl[11509], bl[11510], bl[11511], bl[11512], bl[11513], bl[11514], bl[11515], bl[11516], bl[11517], bl[11518], bl[11519], bl[11520], bl[11521], bl[11522], bl[11523]}),
        .wl({wl[10424], wl[10425], wl[10426], wl[10427], wl[10428], wl[10429], wl[10430], wl[10431], wl[10432], wl[10433], wl[10434], wl[10435], wl[10436], wl[10437], wl[10438], wl[10439], wl[10440], wl[10441], wl[10442], wl[10443], wl[10444], wl[10445], wl[10446], wl[10447], wl[10448], wl[10449], wl[10450], wl[10451], wl[10452], wl[10453], wl[10454], wl[10455], wl[10456], wl[10457], wl[10458], wl[10459], wl[10460], wl[10461], wl[10462], wl[10463], wl[10464], wl[10465], wl[10466], wl[10467], wl[10468], wl[10469], wl[10470], wl[10471], wl[10472], wl[10473], wl[10474], wl[10475], wl[10476], wl[10477], wl[10478], wl[10479], wl[10480], wl[10481], wl[10482], wl[10483], wl[10484], wl[10485], wl[10486], wl[10487], wl[10488], wl[10489], wl[10490], wl[10491], wl[10492], wl[10493], wl[10494], wl[10495], wl[10496], wl[10497], wl[10498], wl[10499], wl[10500], wl[10501], wl[10502], wl[10503], wl[10504], wl[10505], wl[10506], wl[10507], wl[10508], wl[10509], wl[10510], wl[10511], wl[10512], wl[10513], wl[10514], wl[10515], wl[10516], wl[10517], wl[10518], wl[10519], wl[10520], wl[10521], wl[10522], wl[10523], wl[10524], wl[10525], wl[10526], wl[10527], wl[10528], wl[10529], wl[10530], wl[10531], wl[10532], wl[10533], wl[10534], wl[10535], wl[10536], wl[10537], wl[10538], wl[10539], wl[10540], wl[10541], wl[10542], wl[10543], wl[10544], wl[10545], wl[10546], wl[10547], wl[10548], wl[10549], wl[10550], wl[10551], wl[10552], wl[10553], wl[10554], wl[10555], wl[10556], wl[10557], wl[10558], wl[10559], wl[10560], wl[10561], wl[10562], wl[10563], wl[10564], wl[10565], wl[10566], wl[10567], wl[10568], wl[10569], wl[10570], wl[10571], wl[10572], wl[10573], wl[10574], wl[10575], wl[10576], wl[10577], wl[10578], wl[10579], wl[10580], wl[10581], wl[10582], wl[10583], wl[10584], wl[10585], wl[10586], wl[10587], wl[10588], wl[10589], wl[10590], wl[10591], wl[10592], wl[10593], wl[10594], wl[10595], wl[10596], wl[10597], wl[10598], wl[10599], wl[10600], wl[10601], wl[10602], wl[10603], wl[10604], wl[10605], wl[10606], wl[10607], wl[10608], wl[10609], wl[10610], wl[10611], wl[10612], wl[10613], wl[10614], wl[10615], wl[10616], wl[10617], wl[10618], wl[10619], wl[10620], wl[10621], wl[10622], wl[10623], wl[10624], wl[10625], wl[10626], wl[10627], wl[10628], wl[10629], wl[10630], wl[10631], wl[10632], wl[10633], wl[10634], wl[10635], wl[10636], wl[10637], wl[10638], wl[10639], wl[10640], wl[10641], wl[10642], wl[10643], wl[10644], wl[10645], wl[10646], wl[10647], wl[10648], wl[10649], wl[10650], wl[10651], wl[10652], wl[10653], wl[10654], wl[10655], wl[10656], wl[10657], wl[10658], wl[10659], wl[10660], wl[10661], wl[10662], wl[10663], wl[10664], wl[10665], wl[10666], wl[10667], wl[10668], wl[10669], wl[10670], wl[10671], wl[10672], wl[10673], wl[10674], wl[10675], wl[10676], wl[10677], wl[10678], wl[10679], wl[10680], wl[10681], wl[10682], wl[10683], wl[10684], wl[10685], wl[10686], wl[10687], wl[10688], wl[10689], wl[10690], wl[10691], wl[10692], wl[10693], wl[10694], wl[10695], wl[10696], wl[10697], wl[10698], wl[10699], wl[10700], wl[10701], wl[10702], wl[10703], wl[10704], wl[10705], wl[10706], wl[10707], wl[10708], wl[10709], wl[10710], wl[10711], wl[10712], wl[10713], wl[10714], wl[10715], wl[10716], wl[10717], wl[10718], wl[10719], wl[10720], wl[10721], wl[10722], wl[10723], wl[10724], wl[10725], wl[10726], wl[10727], wl[10728], wl[10729], wl[10730], wl[10731], wl[10732], wl[10733], wl[10734], wl[10735], wl[10736], wl[10737], wl[10738], wl[10739], wl[10740], wl[10741], wl[10742], wl[10743], wl[10744], wl[10745], wl[10746], wl[10747], wl[10748], wl[10749], wl[10750], wl[10751], wl[10752], wl[10753], wl[10754], wl[10755], wl[10756], wl[10757], wl[10758], wl[10759], wl[10760], wl[10761], wl[10762], wl[10763], wl[10764], wl[10765], wl[10766], wl[10767], wl[10768], wl[10769], wl[10770], wl[10771], wl[10772], wl[10773], wl[10774], wl[10775], wl[10776], wl[10777], wl[10778], wl[10779], wl[10780], wl[10781], wl[10782], wl[10783], wl[10784], wl[10785], wl[10786], wl[10787], wl[10788], wl[10789], wl[10790], wl[10791], wl[10792], wl[10793], wl[10794], wl[10795], wl[10796], wl[10797], wl[10798], wl[10799], wl[10800], wl[10801], wl[10802], wl[10803], wl[10804], wl[10805], wl[10806], wl[10807], wl[10808], wl[10809], wl[10810], wl[10811], wl[10812], wl[10813], wl[10814], wl[10815], wl[10816], wl[10817], wl[10818], wl[10819], wl[10820], wl[10821], wl[10822], wl[10823], wl[10824], wl[10825], wl[10826], wl[10827], wl[10828], wl[10829], wl[10830], wl[10831], wl[10832], wl[10833], wl[10834], wl[10835], wl[10836], wl[10837], wl[10838], wl[10839], wl[10840], wl[10841], wl[10842], wl[10843], wl[10844], wl[10845], wl[10846], wl[10847], wl[10848], wl[10849], wl[10850], wl[10851], wl[10852], wl[10853], wl[10854], wl[10855], wl[10856], wl[10857], wl[10858], wl[10859], wl[10860], wl[10861], wl[10862], wl[10863], wl[10864], wl[10865], wl[10866], wl[10867], wl[10868], wl[10869], wl[10870], wl[10871], wl[10872], wl[10873], wl[10874], wl[10875], wl[10876], wl[10877], wl[10878], wl[10879], wl[10880], wl[10881], wl[10882], wl[10883], wl[10884], wl[10885], wl[10886], wl[10887], wl[10888], wl[10889], wl[10890], wl[10891], wl[10892], wl[10893], wl[10894], wl[10895], wl[10896], wl[10897], wl[10898], wl[10899], wl[10900], wl[10901], wl[10902], wl[10903], wl[10904], wl[10905], wl[10906], wl[10907], wl[10908], wl[10909], wl[10910], wl[10911], wl[10912], wl[10913], wl[10914], wl[10915], wl[10916], wl[10917], wl[10918], wl[10919], wl[10920], wl[10921], wl[10922], wl[10923], wl[10924], wl[10925], wl[10926], wl[10927], wl[10928], wl[10929], wl[10930], wl[10931], wl[10932], wl[10933], wl[10934], wl[10935], wl[10936], wl[10937], wl[10938], wl[10939], wl[10940], wl[10941], wl[10942], wl[10943], wl[10944], wl[10945], wl[10946], wl[10947], wl[10948], wl[10949], wl[10950], wl[10951], wl[10952], wl[10953], wl[10954], wl[10955], wl[10956], wl[10957], wl[10958], wl[10959], wl[10960], wl[10961], wl[10962], wl[10963], wl[10964], wl[10965], wl[10966], wl[10967], wl[10968], wl[10969], wl[10970], wl[10971], wl[10972], wl[10973], wl[10974], wl[10975], wl[10976], wl[10977], wl[10978], wl[10979], wl[10980], wl[10981], wl[10982], wl[10983], wl[10984], wl[10985], wl[10986], wl[10987], wl[10988], wl[10989], wl[10990], wl[10991], wl[10992], wl[10993], wl[10994], wl[10995], wl[10996], wl[10997], wl[10998], wl[10999], wl[11000], wl[11001], wl[11002], wl[11003], wl[11004], wl[11005], wl[11006], wl[11007], wl[11008], wl[11009], wl[11010], wl[11011], wl[11012], wl[11013], wl[11014], wl[11015], wl[11016], wl[11017], wl[11018], wl[11019], wl[11020], wl[11021], wl[11022], wl[11023], wl[11024], wl[11025], wl[11026], wl[11027], wl[11028], wl[11029], wl[11030], wl[11031], wl[11032], wl[11033], wl[11034], wl[11035], wl[11036], wl[11037], wl[11038], wl[11039], wl[11040], wl[11041], wl[11042], wl[11043], wl[11044], wl[11045], wl[11046], wl[11047], wl[11048], wl[11049], wl[11050], wl[11051], wl[11052], wl[11053], wl[11054], wl[11055], wl[11056], wl[11057], wl[11058], wl[11059], wl[11060], wl[11061], wl[11062], wl[11063], wl[11064], wl[11065], wl[11066], wl[11067], wl[11068], wl[11069], wl[11070], wl[11071], wl[11072], wl[11073], wl[11074], wl[11075], wl[11076], wl[11077], wl[11078], wl[11079], wl[11080], wl[11081], wl[11082], wl[11083], wl[11084], wl[11085], wl[11086], wl[11087], wl[11088], wl[11089], wl[11090], wl[11091], wl[11092], wl[11093], wl[11094], wl[11095], wl[11096], wl[11097], wl[11098], wl[11099], wl[11100], wl[11101], wl[11102], wl[11103], wl[11104], wl[11105], wl[11106], wl[11107], wl[11108], wl[11109], wl[11110], wl[11111], wl[11112], wl[11113], wl[11114], wl[11115], wl[11116], wl[11117], wl[11118], wl[11119], wl[11120], wl[11121], wl[11122], wl[11123], wl[11124], wl[11125], wl[11126], wl[11127], wl[11128], wl[11129], wl[11130], wl[11131], wl[11132], wl[11133], wl[11134], wl[11135], wl[11136], wl[11137], wl[11138], wl[11139], wl[11140], wl[11141], wl[11142], wl[11143], wl[11144], wl[11145], wl[11146], wl[11147], wl[11148], wl[11149], wl[11150], wl[11151], wl[11152], wl[11153], wl[11154], wl[11155], wl[11156], wl[11157], wl[11158], wl[11159], wl[11160], wl[11161], wl[11162], wl[11163], wl[11164], wl[11165], wl[11166], wl[11167], wl[11168], wl[11169], wl[11170], wl[11171], wl[11172], wl[11173], wl[11174], wl[11175], wl[11176], wl[11177], wl[11178], wl[11179], wl[11180], wl[11181], wl[11182], wl[11183], wl[11184], wl[11185], wl[11186], wl[11187], wl[11188], wl[11189], wl[11190], wl[11191], wl[11192], wl[11193], wl[11194], wl[11195], wl[11196], wl[11197], wl[11198], wl[11199], wl[11200], wl[11201], wl[11202], wl[11203], wl[11204], wl[11205], wl[11206], wl[11207], wl[11208], wl[11209], wl[11210], wl[11211], wl[11212], wl[11213], wl[11214], wl[11215], wl[11216], wl[11217], wl[11218], wl[11219], wl[11220], wl[11221], wl[11222], wl[11223], wl[11224], wl[11225], wl[11226], wl[11227], wl[11228], wl[11229], wl[11230], wl[11231], wl[11232], wl[11233], wl[11234], wl[11235], wl[11236], wl[11237], wl[11238], wl[11239], wl[11240], wl[11241], wl[11242], wl[11243], wl[11244], wl[11245], wl[11246], wl[11247], wl[11248], wl[11249], wl[11250], wl[11251], wl[11252], wl[11253], wl[11254], wl[11255], wl[11256], wl[11257], wl[11258], wl[11259], wl[11260], wl[11261], wl[11262], wl[11263], wl[11264], wl[11265], wl[11266], wl[11267], wl[11268], wl[11269], wl[11270], wl[11271], wl[11272], wl[11273], wl[11274], wl[11275], wl[11276], wl[11277], wl[11278], wl[11279], wl[11280], wl[11281], wl[11282], wl[11283], wl[11284], wl[11285], wl[11286], wl[11287], wl[11288], wl[11289], wl[11290], wl[11291], wl[11292], wl[11293], wl[11294], wl[11295], wl[11296], wl[11297], wl[11298], wl[11299], wl[11300], wl[11301], wl[11302], wl[11303], wl[11304], wl[11305], wl[11306], wl[11307], wl[11308], wl[11309], wl[11310], wl[11311], wl[11312], wl[11313], wl[11314], wl[11315], wl[11316], wl[11317], wl[11318], wl[11319], wl[11320], wl[11321], wl[11322], wl[11323], wl[11324], wl[11325], wl[11326], wl[11327], wl[11328], wl[11329], wl[11330], wl[11331], wl[11332], wl[11333], wl[11334], wl[11335], wl[11336], wl[11337], wl[11338], wl[11339], wl[11340], wl[11341], wl[11342], wl[11343], wl[11344], wl[11345], wl[11346], wl[11347], wl[11348], wl[11349], wl[11350], wl[11351], wl[11352], wl[11353], wl[11354], wl[11355], wl[11356], wl[11357], wl[11358], wl[11359], wl[11360], wl[11361], wl[11362], wl[11363], wl[11364], wl[11365], wl[11366], wl[11367], wl[11368], wl[11369], wl[11370], wl[11371], wl[11372], wl[11373], wl[11374], wl[11375], wl[11376], wl[11377], wl[11378], wl[11379], wl[11380], wl[11381], wl[11382], wl[11383], wl[11384], wl[11385], wl[11386], wl[11387], wl[11388], wl[11389], wl[11390], wl[11391], wl[11392], wl[11393], wl[11394], wl[11395], wl[11396], wl[11397], wl[11398], wl[11399], wl[11400], wl[11401], wl[11402], wl[11403], wl[11404], wl[11405], wl[11406], wl[11407], wl[11408], wl[11409], wl[11410], wl[11411], wl[11412], wl[11413], wl[11414], wl[11415], wl[11416], wl[11417], wl[11418], wl[11419], wl[11420], wl[11421], wl[11422], wl[11423], wl[11424], wl[11425], wl[11426], wl[11427], wl[11428], wl[11429], wl[11430], wl[11431], wl[11432], wl[11433], wl[11434], wl[11435], wl[11436], wl[11437], wl[11438], wl[11439], wl[11440], wl[11441], wl[11442], wl[11443], wl[11524], wl[11525], wl[11526], wl[11527], wl[11528], wl[11529], wl[11530], wl[11531], wl[11532], wl[11533], wl[11534], wl[11535], wl[11536], wl[11537], wl[11538], wl[11539], wl[11540], wl[11541], wl[11542], wl[11543], wl[11544], wl[11545], wl[11546], wl[11547], wl[11548], wl[11549], wl[11550], wl[11551], wl[11552], wl[11553], wl[11554], wl[11555], wl[11556], wl[11557], wl[11558], wl[11559], wl[11560], wl[11561], wl[11562], wl[11563], wl[11564], wl[11565], wl[11566], wl[11567], wl[11568], wl[11569], wl[11570], wl[11571], wl[11572], wl[11573], wl[11574], wl[11575], wl[11576], wl[11577], wl[11578], wl[11579], wl[11580], wl[11581], wl[11582], wl[11583], wl[11584], wl[11585], wl[11586], wl[11587], wl[11588], wl[11589], wl[11590], wl[11591], wl[11592], wl[11593], wl[11594], wl[11595], wl[11596], wl[11597], wl[11598], wl[11599], wl[11600], wl[11601], wl[11602], wl[11603], wl[10344], wl[10345], wl[10346], wl[10347], wl[10348], wl[10349], wl[10350], wl[10351], wl[10352], wl[10353], wl[10354], wl[10355], wl[10356], wl[10357], wl[10358], wl[10359], wl[10360], wl[10361], wl[10362], wl[10363], wl[10364], wl[10365], wl[10366], wl[10367], wl[10368], wl[10369], wl[10370], wl[10371], wl[10372], wl[10373], wl[10374], wl[10375], wl[10376], wl[10377], wl[10378], wl[10379], wl[10380], wl[10381], wl[10382], wl[10383], wl[10384], wl[10385], wl[10386], wl[10387], wl[10388], wl[10389], wl[10390], wl[10391], wl[10392], wl[10393], wl[10394], wl[10395], wl[10396], wl[10397], wl[10398], wl[10399], wl[10400], wl[10401], wl[10402], wl[10403], wl[10404], wl[10405], wl[10406], wl[10407], wl[10408], wl[10409], wl[10410], wl[10411], wl[10412], wl[10413], wl[10414], wl[10415], wl[10416], wl[10417], wl[10418], wl[10419], wl[10420], wl[10421], wl[10422], wl[10423], wl[11444], wl[11445], wl[11446], wl[11447], wl[11448], wl[11449], wl[11450], wl[11451], wl[11452], wl[11453], wl[11454], wl[11455], wl[11456], wl[11457], wl[11458], wl[11459], wl[11460], wl[11461], wl[11462], wl[11463], wl[11464], wl[11465], wl[11466], wl[11467], wl[11468], wl[11469], wl[11470], wl[11471], wl[11472], wl[11473], wl[11474], wl[11475], wl[11476], wl[11477], wl[11478], wl[11479], wl[11480], wl[11481], wl[11482], wl[11483], wl[11484], wl[11485], wl[11486], wl[11487], wl[11488], wl[11489], wl[11490], wl[11491], wl[11492], wl[11493], wl[11494], wl[11495], wl[11496], wl[11497], wl[11498], wl[11499], wl[11500], wl[11501], wl[11502], wl[11503], wl[11504], wl[11505], wl[11506], wl[11507], wl[11508], wl[11509], wl[11510], wl[11511], wl[11512], wl[11513], wl[11514], wl[11515], wl[11516], wl[11517], wl[11518], wl[11519], wl[11520], wl[11521], wl[11522], wl[11523]})
    );
    tile tile_2__4_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_0__3__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_0__3__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_0__3__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_1__2__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_1__2__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_1__2__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_0__2__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_0__2__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_0__2__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_0__2__grid_top_r_in[1]),
        .grid_left_in(grid_clb_1__3__grid_left_in),
        .grid_bottom_in(grid_clb_1__3__grid_bottom_in),
        .chanx_left_in(sb_0__1__2_chanx_right_out),
        .chanx_left_out(cbx_1__1__2_chanx_left_out),
        .grid_top_out(grid_clb_1__4__grid_bottom_in),
        .chany_bottom_in(sb_1__1__1_chany_top_out),
        .chany_bottom_out(cby_1__1__2_chany_bottom_out),
        .grid_right_out(grid_clb_2__3__grid_left_in),
        .chany_top_in_0(cby_1__1__3_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__5_chanx_left_out),
        .chany_top_out_0(sb_1__1__2_chany_top_out),
        .chanx_right_out_0(sb_1__1__2_chanx_right_out),
        .grid_top_r_in(sb_1__3__grid_top_r_in),
        .grid_top_l_in(sb_1__3__grid_top_l_in),
        .grid_right_t_in(sb_1__3__grid_right_t_in),
        .grid_right_b_in(sb_1__3__grid_right_b_in),
        .grid_bottom_r_in(sb_1__2__grid_top_r_in),
        .grid_bottom_l_in(sb_1__2__grid_top_l_in),
        .grid_left_t_in(sb_0__3__grid_right_t_in),
        .grid_left_b_in(sb_0__3__grid_right_b_in),
        .bl({bl[11684], bl[11685], bl[11686], bl[11687], bl[11688], bl[11689], bl[11690], bl[11691], bl[11692], bl[11693], bl[11694], bl[11695], bl[11696], bl[11697], bl[11698], bl[11699], bl[11700], bl[11701], bl[11702], bl[11703], bl[11704], bl[11705], bl[11706], bl[11707], bl[11708], bl[11709], bl[11710], bl[11711], bl[11712], bl[11713], bl[11714], bl[11715], bl[11716], bl[11717], bl[11718], bl[11719], bl[11720], bl[11721], bl[11722], bl[11723], bl[11724], bl[11725], bl[11726], bl[11727], bl[11728], bl[11729], bl[11730], bl[11731], bl[11732], bl[11733], bl[11734], bl[11735], bl[11736], bl[11737], bl[11738], bl[11739], bl[11740], bl[11741], bl[11742], bl[11743], bl[11744], bl[11745], bl[11746], bl[11747], bl[11748], bl[11749], bl[11750], bl[11751], bl[11752], bl[11753], bl[11754], bl[11755], bl[11756], bl[11757], bl[11758], bl[11759], bl[11760], bl[11761], bl[11762], bl[11763], bl[11764], bl[11765], bl[11766], bl[11767], bl[11768], bl[11769], bl[11770], bl[11771], bl[11772], bl[11773], bl[11774], bl[11775], bl[11776], bl[11777], bl[11778], bl[11779], bl[11780], bl[11781], bl[11782], bl[11783], bl[11784], bl[11785], bl[11786], bl[11787], bl[11788], bl[11789], bl[11790], bl[11791], bl[11792], bl[11793], bl[11794], bl[11795], bl[11796], bl[11797], bl[11798], bl[11799], bl[11800], bl[11801], bl[11802], bl[11803], bl[11804], bl[11805], bl[11806], bl[11807], bl[11808], bl[11809], bl[11810], bl[11811], bl[11812], bl[11813], bl[11814], bl[11815], bl[11816], bl[11817], bl[11818], bl[11819], bl[11820], bl[11821], bl[11822], bl[11823], bl[11824], bl[11825], bl[11826], bl[11827], bl[11828], bl[11829], bl[11830], bl[11831], bl[11832], bl[11833], bl[11834], bl[11835], bl[11836], bl[11837], bl[11838], bl[11839], bl[11840], bl[11841], bl[11842], bl[11843], bl[11844], bl[11845], bl[11846], bl[11847], bl[11848], bl[11849], bl[11850], bl[11851], bl[11852], bl[11853], bl[11854], bl[11855], bl[11856], bl[11857], bl[11858], bl[11859], bl[11860], bl[11861], bl[11862], bl[11863], bl[11864], bl[11865], bl[11866], bl[11867], bl[11868], bl[11869], bl[11870], bl[11871], bl[11872], bl[11873], bl[11874], bl[11875], bl[11876], bl[11877], bl[11878], bl[11879], bl[11880], bl[11881], bl[11882], bl[11883], bl[11884], bl[11885], bl[11886], bl[11887], bl[11888], bl[11889], bl[11890], bl[11891], bl[11892], bl[11893], bl[11894], bl[11895], bl[11896], bl[11897], bl[11898], bl[11899], bl[11900], bl[11901], bl[11902], bl[11903], bl[11904], bl[11905], bl[11906], bl[11907], bl[11908], bl[11909], bl[11910], bl[11911], bl[11912], bl[11913], bl[11914], bl[11915], bl[11916], bl[11917], bl[11918], bl[11919], bl[11920], bl[11921], bl[11922], bl[11923], bl[11924], bl[11925], bl[11926], bl[11927], bl[11928], bl[11929], bl[11930], bl[11931], bl[11932], bl[11933], bl[11934], bl[11935], bl[11936], bl[11937], bl[11938], bl[11939], bl[11940], bl[11941], bl[11942], bl[11943], bl[11944], bl[11945], bl[11946], bl[11947], bl[11948], bl[11949], bl[11950], bl[11951], bl[11952], bl[11953], bl[11954], bl[11955], bl[11956], bl[11957], bl[11958], bl[11959], bl[11960], bl[11961], bl[11962], bl[11963], bl[11964], bl[11965], bl[11966], bl[11967], bl[11968], bl[11969], bl[11970], bl[11971], bl[11972], bl[11973], bl[11974], bl[11975], bl[11976], bl[11977], bl[11978], bl[11979], bl[11980], bl[11981], bl[11982], bl[11983], bl[11984], bl[11985], bl[11986], bl[11987], bl[11988], bl[11989], bl[11990], bl[11991], bl[11992], bl[11993], bl[11994], bl[11995], bl[11996], bl[11997], bl[11998], bl[11999], bl[12000], bl[12001], bl[12002], bl[12003], bl[12004], bl[12005], bl[12006], bl[12007], bl[12008], bl[12009], bl[12010], bl[12011], bl[12012], bl[12013], bl[12014], bl[12015], bl[12016], bl[12017], bl[12018], bl[12019], bl[12020], bl[12021], bl[12022], bl[12023], bl[12024], bl[12025], bl[12026], bl[12027], bl[12028], bl[12029], bl[12030], bl[12031], bl[12032], bl[12033], bl[12034], bl[12035], bl[12036], bl[12037], bl[12038], bl[12039], bl[12040], bl[12041], bl[12042], bl[12043], bl[12044], bl[12045], bl[12046], bl[12047], bl[12048], bl[12049], bl[12050], bl[12051], bl[12052], bl[12053], bl[12054], bl[12055], bl[12056], bl[12057], bl[12058], bl[12059], bl[12060], bl[12061], bl[12062], bl[12063], bl[12064], bl[12065], bl[12066], bl[12067], bl[12068], bl[12069], bl[12070], bl[12071], bl[12072], bl[12073], bl[12074], bl[12075], bl[12076], bl[12077], bl[12078], bl[12079], bl[12080], bl[12081], bl[12082], bl[12083], bl[12084], bl[12085], bl[12086], bl[12087], bl[12088], bl[12089], bl[12090], bl[12091], bl[12092], bl[12093], bl[12094], bl[12095], bl[12096], bl[12097], bl[12098], bl[12099], bl[12100], bl[12101], bl[12102], bl[12103], bl[12104], bl[12105], bl[12106], bl[12107], bl[12108], bl[12109], bl[12110], bl[12111], bl[12112], bl[12113], bl[12114], bl[12115], bl[12116], bl[12117], bl[12118], bl[12119], bl[12120], bl[12121], bl[12122], bl[12123], bl[12124], bl[12125], bl[12126], bl[12127], bl[12128], bl[12129], bl[12130], bl[12131], bl[12132], bl[12133], bl[12134], bl[12135], bl[12136], bl[12137], bl[12138], bl[12139], bl[12140], bl[12141], bl[12142], bl[12143], bl[12144], bl[12145], bl[12146], bl[12147], bl[12148], bl[12149], bl[12150], bl[12151], bl[12152], bl[12153], bl[12154], bl[12155], bl[12156], bl[12157], bl[12158], bl[12159], bl[12160], bl[12161], bl[12162], bl[12163], bl[12164], bl[12165], bl[12166], bl[12167], bl[12168], bl[12169], bl[12170], bl[12171], bl[12172], bl[12173], bl[12174], bl[12175], bl[12176], bl[12177], bl[12178], bl[12179], bl[12180], bl[12181], bl[12182], bl[12183], bl[12184], bl[12185], bl[12186], bl[12187], bl[12188], bl[12189], bl[12190], bl[12191], bl[12192], bl[12193], bl[12194], bl[12195], bl[12196], bl[12197], bl[12198], bl[12199], bl[12200], bl[12201], bl[12202], bl[12203], bl[12204], bl[12205], bl[12206], bl[12207], bl[12208], bl[12209], bl[12210], bl[12211], bl[12212], bl[12213], bl[12214], bl[12215], bl[12216], bl[12217], bl[12218], bl[12219], bl[12220], bl[12221], bl[12222], bl[12223], bl[12224], bl[12225], bl[12226], bl[12227], bl[12228], bl[12229], bl[12230], bl[12231], bl[12232], bl[12233], bl[12234], bl[12235], bl[12236], bl[12237], bl[12238], bl[12239], bl[12240], bl[12241], bl[12242], bl[12243], bl[12244], bl[12245], bl[12246], bl[12247], bl[12248], bl[12249], bl[12250], bl[12251], bl[12252], bl[12253], bl[12254], bl[12255], bl[12256], bl[12257], bl[12258], bl[12259], bl[12260], bl[12261], bl[12262], bl[12263], bl[12264], bl[12265], bl[12266], bl[12267], bl[12268], bl[12269], bl[12270], bl[12271], bl[12272], bl[12273], bl[12274], bl[12275], bl[12276], bl[12277], bl[12278], bl[12279], bl[12280], bl[12281], bl[12282], bl[12283], bl[12284], bl[12285], bl[12286], bl[12287], bl[12288], bl[12289], bl[12290], bl[12291], bl[12292], bl[12293], bl[12294], bl[12295], bl[12296], bl[12297], bl[12298], bl[12299], bl[12300], bl[12301], bl[12302], bl[12303], bl[12304], bl[12305], bl[12306], bl[12307], bl[12308], bl[12309], bl[12310], bl[12311], bl[12312], bl[12313], bl[12314], bl[12315], bl[12316], bl[12317], bl[12318], bl[12319], bl[12320], bl[12321], bl[12322], bl[12323], bl[12324], bl[12325], bl[12326], bl[12327], bl[12328], bl[12329], bl[12330], bl[12331], bl[12332], bl[12333], bl[12334], bl[12335], bl[12336], bl[12337], bl[12338], bl[12339], bl[12340], bl[12341], bl[12342], bl[12343], bl[12344], bl[12345], bl[12346], bl[12347], bl[12348], bl[12349], bl[12350], bl[12351], bl[12352], bl[12353], bl[12354], bl[12355], bl[12356], bl[12357], bl[12358], bl[12359], bl[12360], bl[12361], bl[12362], bl[12363], bl[12364], bl[12365], bl[12366], bl[12367], bl[12368], bl[12369], bl[12370], bl[12371], bl[12372], bl[12373], bl[12374], bl[12375], bl[12376], bl[12377], bl[12378], bl[12379], bl[12380], bl[12381], bl[12382], bl[12383], bl[12384], bl[12385], bl[12386], bl[12387], bl[12388], bl[12389], bl[12390], bl[12391], bl[12392], bl[12393], bl[12394], bl[12395], bl[12396], bl[12397], bl[12398], bl[12399], bl[12400], bl[12401], bl[12402], bl[12403], bl[12404], bl[12405], bl[12406], bl[12407], bl[12408], bl[12409], bl[12410], bl[12411], bl[12412], bl[12413], bl[12414], bl[12415], bl[12416], bl[12417], bl[12418], bl[12419], bl[12420], bl[12421], bl[12422], bl[12423], bl[12424], bl[12425], bl[12426], bl[12427], bl[12428], bl[12429], bl[12430], bl[12431], bl[12432], bl[12433], bl[12434], bl[12435], bl[12436], bl[12437], bl[12438], bl[12439], bl[12440], bl[12441], bl[12442], bl[12443], bl[12444], bl[12445], bl[12446], bl[12447], bl[12448], bl[12449], bl[12450], bl[12451], bl[12452], bl[12453], bl[12454], bl[12455], bl[12456], bl[12457], bl[12458], bl[12459], bl[12460], bl[12461], bl[12462], bl[12463], bl[12464], bl[12465], bl[12466], bl[12467], bl[12468], bl[12469], bl[12470], bl[12471], bl[12472], bl[12473], bl[12474], bl[12475], bl[12476], bl[12477], bl[12478], bl[12479], bl[12480], bl[12481], bl[12482], bl[12483], bl[12484], bl[12485], bl[12486], bl[12487], bl[12488], bl[12489], bl[12490], bl[12491], bl[12492], bl[12493], bl[12494], bl[12495], bl[12496], bl[12497], bl[12498], bl[12499], bl[12500], bl[12501], bl[12502], bl[12503], bl[12504], bl[12505], bl[12506], bl[12507], bl[12508], bl[12509], bl[12510], bl[12511], bl[12512], bl[12513], bl[12514], bl[12515], bl[12516], bl[12517], bl[12518], bl[12519], bl[12520], bl[12521], bl[12522], bl[12523], bl[12524], bl[12525], bl[12526], bl[12527], bl[12528], bl[12529], bl[12530], bl[12531], bl[12532], bl[12533], bl[12534], bl[12535], bl[12536], bl[12537], bl[12538], bl[12539], bl[12540], bl[12541], bl[12542], bl[12543], bl[12544], bl[12545], bl[12546], bl[12547], bl[12548], bl[12549], bl[12550], bl[12551], bl[12552], bl[12553], bl[12554], bl[12555], bl[12556], bl[12557], bl[12558], bl[12559], bl[12560], bl[12561], bl[12562], bl[12563], bl[12564], bl[12565], bl[12566], bl[12567], bl[12568], bl[12569], bl[12570], bl[12571], bl[12572], bl[12573], bl[12574], bl[12575], bl[12576], bl[12577], bl[12578], bl[12579], bl[12580], bl[12581], bl[12582], bl[12583], bl[12584], bl[12585], bl[12586], bl[12587], bl[12588], bl[12589], bl[12590], bl[12591], bl[12592], bl[12593], bl[12594], bl[12595], bl[12596], bl[12597], bl[12598], bl[12599], bl[12600], bl[12601], bl[12602], bl[12603], bl[12604], bl[12605], bl[12606], bl[12607], bl[12608], bl[12609], bl[12610], bl[12611], bl[12612], bl[12613], bl[12614], bl[12615], bl[12616], bl[12617], bl[12618], bl[12619], bl[12620], bl[12621], bl[12622], bl[12623], bl[12624], bl[12625], bl[12626], bl[12627], bl[12628], bl[12629], bl[12630], bl[12631], bl[12632], bl[12633], bl[12634], bl[12635], bl[12636], bl[12637], bl[12638], bl[12639], bl[12640], bl[12641], bl[12642], bl[12643], bl[12644], bl[12645], bl[12646], bl[12647], bl[12648], bl[12649], bl[12650], bl[12651], bl[12652], bl[12653], bl[12654], bl[12655], bl[12656], bl[12657], bl[12658], bl[12659], bl[12660], bl[12661], bl[12662], bl[12663], bl[12664], bl[12665], bl[12666], bl[12667], bl[12668], bl[12669], bl[12670], bl[12671], bl[12672], bl[12673], bl[12674], bl[12675], bl[12676], bl[12677], bl[12678], bl[12679], bl[12680], bl[12681], bl[12682], bl[12683], bl[12684], bl[12685], bl[12686], bl[12687], bl[12688], bl[12689], bl[12690], bl[12691], bl[12692], bl[12693], bl[12694], bl[12695], bl[12696], bl[12697], bl[12698], bl[12699], bl[12700], bl[12701], bl[12702], bl[12703], bl[20328], bl[20329], bl[20330], bl[20331], bl[20332], bl[20333], bl[20334], bl[20335], bl[20336], bl[20337], bl[20338], bl[20339], bl[20340], bl[20341], bl[20342], bl[20343], bl[20344], bl[20345], bl[20346], bl[20347], bl[20348], bl[20349], bl[20350], bl[20351], bl[20352], bl[20353], bl[20354], bl[20355], bl[20356], bl[20357], bl[20358], bl[20359], bl[20360], bl[20361], bl[20362], bl[20363], bl[20364], bl[20365], bl[20366], bl[20367], bl[20368], bl[20369], bl[20370], bl[20371], bl[20372], bl[20373], bl[20374], bl[20375], bl[20376], bl[20377], bl[20378], bl[20379], bl[20380], bl[20381], bl[20382], bl[20383], bl[20384], bl[20385], bl[20386], bl[20387], bl[20388], bl[20389], bl[20390], bl[20391], bl[20392], bl[20393], bl[20394], bl[20395], bl[20396], bl[20397], bl[20398], bl[20399], bl[20400], bl[20401], bl[20402], bl[20403], bl[20404], bl[20405], bl[20406], bl[20407], bl[11604], bl[11605], bl[11606], bl[11607], bl[11608], bl[11609], bl[11610], bl[11611], bl[11612], bl[11613], bl[11614], bl[11615], bl[11616], bl[11617], bl[11618], bl[11619], bl[11620], bl[11621], bl[11622], bl[11623], bl[11624], bl[11625], bl[11626], bl[11627], bl[11628], bl[11629], bl[11630], bl[11631], bl[11632], bl[11633], bl[11634], bl[11635], bl[11636], bl[11637], bl[11638], bl[11639], bl[11640], bl[11641], bl[11642], bl[11643], bl[11644], bl[11645], bl[11646], bl[11647], bl[11648], bl[11649], bl[11650], bl[11651], bl[11652], bl[11653], bl[11654], bl[11655], bl[11656], bl[11657], bl[11658], bl[11659], bl[11660], bl[11661], bl[11662], bl[11663], bl[11664], bl[11665], bl[11666], bl[11667], bl[11668], bl[11669], bl[11670], bl[11671], bl[11672], bl[11673], bl[11674], bl[11675], bl[11676], bl[11677], bl[11678], bl[11679], bl[11680], bl[11681], bl[11682], bl[11683], bl[20248], bl[20249], bl[20250], bl[20251], bl[20252], bl[20253], bl[20254], bl[20255], bl[20256], bl[20257], bl[20258], bl[20259], bl[20260], bl[20261], bl[20262], bl[20263], bl[20264], bl[20265], bl[20266], bl[20267], bl[20268], bl[20269], bl[20270], bl[20271], bl[20272], bl[20273], bl[20274], bl[20275], bl[20276], bl[20277], bl[20278], bl[20279], bl[20280], bl[20281], bl[20282], bl[20283], bl[20284], bl[20285], bl[20286], bl[20287], bl[20288], bl[20289], bl[20290], bl[20291], bl[20292], bl[20293], bl[20294], bl[20295], bl[20296], bl[20297], bl[20298], bl[20299], bl[20300], bl[20301], bl[20302], bl[20303], bl[20304], bl[20305], bl[20306], bl[20307], bl[20308], bl[20309], bl[20310], bl[20311], bl[20312], bl[20313], bl[20314], bl[20315], bl[20316], bl[20317], bl[20318], bl[20319], bl[20320], bl[20321], bl[20322], bl[20323], bl[20324], bl[20325], bl[20326], bl[20327]}),
        .wl({wl[11684], wl[11685], wl[11686], wl[11687], wl[11688], wl[11689], wl[11690], wl[11691], wl[11692], wl[11693], wl[11694], wl[11695], wl[11696], wl[11697], wl[11698], wl[11699], wl[11700], wl[11701], wl[11702], wl[11703], wl[11704], wl[11705], wl[11706], wl[11707], wl[11708], wl[11709], wl[11710], wl[11711], wl[11712], wl[11713], wl[11714], wl[11715], wl[11716], wl[11717], wl[11718], wl[11719], wl[11720], wl[11721], wl[11722], wl[11723], wl[11724], wl[11725], wl[11726], wl[11727], wl[11728], wl[11729], wl[11730], wl[11731], wl[11732], wl[11733], wl[11734], wl[11735], wl[11736], wl[11737], wl[11738], wl[11739], wl[11740], wl[11741], wl[11742], wl[11743], wl[11744], wl[11745], wl[11746], wl[11747], wl[11748], wl[11749], wl[11750], wl[11751], wl[11752], wl[11753], wl[11754], wl[11755], wl[11756], wl[11757], wl[11758], wl[11759], wl[11760], wl[11761], wl[11762], wl[11763], wl[11764], wl[11765], wl[11766], wl[11767], wl[11768], wl[11769], wl[11770], wl[11771], wl[11772], wl[11773], wl[11774], wl[11775], wl[11776], wl[11777], wl[11778], wl[11779], wl[11780], wl[11781], wl[11782], wl[11783], wl[11784], wl[11785], wl[11786], wl[11787], wl[11788], wl[11789], wl[11790], wl[11791], wl[11792], wl[11793], wl[11794], wl[11795], wl[11796], wl[11797], wl[11798], wl[11799], wl[11800], wl[11801], wl[11802], wl[11803], wl[11804], wl[11805], wl[11806], wl[11807], wl[11808], wl[11809], wl[11810], wl[11811], wl[11812], wl[11813], wl[11814], wl[11815], wl[11816], wl[11817], wl[11818], wl[11819], wl[11820], wl[11821], wl[11822], wl[11823], wl[11824], wl[11825], wl[11826], wl[11827], wl[11828], wl[11829], wl[11830], wl[11831], wl[11832], wl[11833], wl[11834], wl[11835], wl[11836], wl[11837], wl[11838], wl[11839], wl[11840], wl[11841], wl[11842], wl[11843], wl[11844], wl[11845], wl[11846], wl[11847], wl[11848], wl[11849], wl[11850], wl[11851], wl[11852], wl[11853], wl[11854], wl[11855], wl[11856], wl[11857], wl[11858], wl[11859], wl[11860], wl[11861], wl[11862], wl[11863], wl[11864], wl[11865], wl[11866], wl[11867], wl[11868], wl[11869], wl[11870], wl[11871], wl[11872], wl[11873], wl[11874], wl[11875], wl[11876], wl[11877], wl[11878], wl[11879], wl[11880], wl[11881], wl[11882], wl[11883], wl[11884], wl[11885], wl[11886], wl[11887], wl[11888], wl[11889], wl[11890], wl[11891], wl[11892], wl[11893], wl[11894], wl[11895], wl[11896], wl[11897], wl[11898], wl[11899], wl[11900], wl[11901], wl[11902], wl[11903], wl[11904], wl[11905], wl[11906], wl[11907], wl[11908], wl[11909], wl[11910], wl[11911], wl[11912], wl[11913], wl[11914], wl[11915], wl[11916], wl[11917], wl[11918], wl[11919], wl[11920], wl[11921], wl[11922], wl[11923], wl[11924], wl[11925], wl[11926], wl[11927], wl[11928], wl[11929], wl[11930], wl[11931], wl[11932], wl[11933], wl[11934], wl[11935], wl[11936], wl[11937], wl[11938], wl[11939], wl[11940], wl[11941], wl[11942], wl[11943], wl[11944], wl[11945], wl[11946], wl[11947], wl[11948], wl[11949], wl[11950], wl[11951], wl[11952], wl[11953], wl[11954], wl[11955], wl[11956], wl[11957], wl[11958], wl[11959], wl[11960], wl[11961], wl[11962], wl[11963], wl[11964], wl[11965], wl[11966], wl[11967], wl[11968], wl[11969], wl[11970], wl[11971], wl[11972], wl[11973], wl[11974], wl[11975], wl[11976], wl[11977], wl[11978], wl[11979], wl[11980], wl[11981], wl[11982], wl[11983], wl[11984], wl[11985], wl[11986], wl[11987], wl[11988], wl[11989], wl[11990], wl[11991], wl[11992], wl[11993], wl[11994], wl[11995], wl[11996], wl[11997], wl[11998], wl[11999], wl[12000], wl[12001], wl[12002], wl[12003], wl[12004], wl[12005], wl[12006], wl[12007], wl[12008], wl[12009], wl[12010], wl[12011], wl[12012], wl[12013], wl[12014], wl[12015], wl[12016], wl[12017], wl[12018], wl[12019], wl[12020], wl[12021], wl[12022], wl[12023], wl[12024], wl[12025], wl[12026], wl[12027], wl[12028], wl[12029], wl[12030], wl[12031], wl[12032], wl[12033], wl[12034], wl[12035], wl[12036], wl[12037], wl[12038], wl[12039], wl[12040], wl[12041], wl[12042], wl[12043], wl[12044], wl[12045], wl[12046], wl[12047], wl[12048], wl[12049], wl[12050], wl[12051], wl[12052], wl[12053], wl[12054], wl[12055], wl[12056], wl[12057], wl[12058], wl[12059], wl[12060], wl[12061], wl[12062], wl[12063], wl[12064], wl[12065], wl[12066], wl[12067], wl[12068], wl[12069], wl[12070], wl[12071], wl[12072], wl[12073], wl[12074], wl[12075], wl[12076], wl[12077], wl[12078], wl[12079], wl[12080], wl[12081], wl[12082], wl[12083], wl[12084], wl[12085], wl[12086], wl[12087], wl[12088], wl[12089], wl[12090], wl[12091], wl[12092], wl[12093], wl[12094], wl[12095], wl[12096], wl[12097], wl[12098], wl[12099], wl[12100], wl[12101], wl[12102], wl[12103], wl[12104], wl[12105], wl[12106], wl[12107], wl[12108], wl[12109], wl[12110], wl[12111], wl[12112], wl[12113], wl[12114], wl[12115], wl[12116], wl[12117], wl[12118], wl[12119], wl[12120], wl[12121], wl[12122], wl[12123], wl[12124], wl[12125], wl[12126], wl[12127], wl[12128], wl[12129], wl[12130], wl[12131], wl[12132], wl[12133], wl[12134], wl[12135], wl[12136], wl[12137], wl[12138], wl[12139], wl[12140], wl[12141], wl[12142], wl[12143], wl[12144], wl[12145], wl[12146], wl[12147], wl[12148], wl[12149], wl[12150], wl[12151], wl[12152], wl[12153], wl[12154], wl[12155], wl[12156], wl[12157], wl[12158], wl[12159], wl[12160], wl[12161], wl[12162], wl[12163], wl[12164], wl[12165], wl[12166], wl[12167], wl[12168], wl[12169], wl[12170], wl[12171], wl[12172], wl[12173], wl[12174], wl[12175], wl[12176], wl[12177], wl[12178], wl[12179], wl[12180], wl[12181], wl[12182], wl[12183], wl[12184], wl[12185], wl[12186], wl[12187], wl[12188], wl[12189], wl[12190], wl[12191], wl[12192], wl[12193], wl[12194], wl[12195], wl[12196], wl[12197], wl[12198], wl[12199], wl[12200], wl[12201], wl[12202], wl[12203], wl[12204], wl[12205], wl[12206], wl[12207], wl[12208], wl[12209], wl[12210], wl[12211], wl[12212], wl[12213], wl[12214], wl[12215], wl[12216], wl[12217], wl[12218], wl[12219], wl[12220], wl[12221], wl[12222], wl[12223], wl[12224], wl[12225], wl[12226], wl[12227], wl[12228], wl[12229], wl[12230], wl[12231], wl[12232], wl[12233], wl[12234], wl[12235], wl[12236], wl[12237], wl[12238], wl[12239], wl[12240], wl[12241], wl[12242], wl[12243], wl[12244], wl[12245], wl[12246], wl[12247], wl[12248], wl[12249], wl[12250], wl[12251], wl[12252], wl[12253], wl[12254], wl[12255], wl[12256], wl[12257], wl[12258], wl[12259], wl[12260], wl[12261], wl[12262], wl[12263], wl[12264], wl[12265], wl[12266], wl[12267], wl[12268], wl[12269], wl[12270], wl[12271], wl[12272], wl[12273], wl[12274], wl[12275], wl[12276], wl[12277], wl[12278], wl[12279], wl[12280], wl[12281], wl[12282], wl[12283], wl[12284], wl[12285], wl[12286], wl[12287], wl[12288], wl[12289], wl[12290], wl[12291], wl[12292], wl[12293], wl[12294], wl[12295], wl[12296], wl[12297], wl[12298], wl[12299], wl[12300], wl[12301], wl[12302], wl[12303], wl[12304], wl[12305], wl[12306], wl[12307], wl[12308], wl[12309], wl[12310], wl[12311], wl[12312], wl[12313], wl[12314], wl[12315], wl[12316], wl[12317], wl[12318], wl[12319], wl[12320], wl[12321], wl[12322], wl[12323], wl[12324], wl[12325], wl[12326], wl[12327], wl[12328], wl[12329], wl[12330], wl[12331], wl[12332], wl[12333], wl[12334], wl[12335], wl[12336], wl[12337], wl[12338], wl[12339], wl[12340], wl[12341], wl[12342], wl[12343], wl[12344], wl[12345], wl[12346], wl[12347], wl[12348], wl[12349], wl[12350], wl[12351], wl[12352], wl[12353], wl[12354], wl[12355], wl[12356], wl[12357], wl[12358], wl[12359], wl[12360], wl[12361], wl[12362], wl[12363], wl[12364], wl[12365], wl[12366], wl[12367], wl[12368], wl[12369], wl[12370], wl[12371], wl[12372], wl[12373], wl[12374], wl[12375], wl[12376], wl[12377], wl[12378], wl[12379], wl[12380], wl[12381], wl[12382], wl[12383], wl[12384], wl[12385], wl[12386], wl[12387], wl[12388], wl[12389], wl[12390], wl[12391], wl[12392], wl[12393], wl[12394], wl[12395], wl[12396], wl[12397], wl[12398], wl[12399], wl[12400], wl[12401], wl[12402], wl[12403], wl[12404], wl[12405], wl[12406], wl[12407], wl[12408], wl[12409], wl[12410], wl[12411], wl[12412], wl[12413], wl[12414], wl[12415], wl[12416], wl[12417], wl[12418], wl[12419], wl[12420], wl[12421], wl[12422], wl[12423], wl[12424], wl[12425], wl[12426], wl[12427], wl[12428], wl[12429], wl[12430], wl[12431], wl[12432], wl[12433], wl[12434], wl[12435], wl[12436], wl[12437], wl[12438], wl[12439], wl[12440], wl[12441], wl[12442], wl[12443], wl[12444], wl[12445], wl[12446], wl[12447], wl[12448], wl[12449], wl[12450], wl[12451], wl[12452], wl[12453], wl[12454], wl[12455], wl[12456], wl[12457], wl[12458], wl[12459], wl[12460], wl[12461], wl[12462], wl[12463], wl[12464], wl[12465], wl[12466], wl[12467], wl[12468], wl[12469], wl[12470], wl[12471], wl[12472], wl[12473], wl[12474], wl[12475], wl[12476], wl[12477], wl[12478], wl[12479], wl[12480], wl[12481], wl[12482], wl[12483], wl[12484], wl[12485], wl[12486], wl[12487], wl[12488], wl[12489], wl[12490], wl[12491], wl[12492], wl[12493], wl[12494], wl[12495], wl[12496], wl[12497], wl[12498], wl[12499], wl[12500], wl[12501], wl[12502], wl[12503], wl[12504], wl[12505], wl[12506], wl[12507], wl[12508], wl[12509], wl[12510], wl[12511], wl[12512], wl[12513], wl[12514], wl[12515], wl[12516], wl[12517], wl[12518], wl[12519], wl[12520], wl[12521], wl[12522], wl[12523], wl[12524], wl[12525], wl[12526], wl[12527], wl[12528], wl[12529], wl[12530], wl[12531], wl[12532], wl[12533], wl[12534], wl[12535], wl[12536], wl[12537], wl[12538], wl[12539], wl[12540], wl[12541], wl[12542], wl[12543], wl[12544], wl[12545], wl[12546], wl[12547], wl[12548], wl[12549], wl[12550], wl[12551], wl[12552], wl[12553], wl[12554], wl[12555], wl[12556], wl[12557], wl[12558], wl[12559], wl[12560], wl[12561], wl[12562], wl[12563], wl[12564], wl[12565], wl[12566], wl[12567], wl[12568], wl[12569], wl[12570], wl[12571], wl[12572], wl[12573], wl[12574], wl[12575], wl[12576], wl[12577], wl[12578], wl[12579], wl[12580], wl[12581], wl[12582], wl[12583], wl[12584], wl[12585], wl[12586], wl[12587], wl[12588], wl[12589], wl[12590], wl[12591], wl[12592], wl[12593], wl[12594], wl[12595], wl[12596], wl[12597], wl[12598], wl[12599], wl[12600], wl[12601], wl[12602], wl[12603], wl[12604], wl[12605], wl[12606], wl[12607], wl[12608], wl[12609], wl[12610], wl[12611], wl[12612], wl[12613], wl[12614], wl[12615], wl[12616], wl[12617], wl[12618], wl[12619], wl[12620], wl[12621], wl[12622], wl[12623], wl[12624], wl[12625], wl[12626], wl[12627], wl[12628], wl[12629], wl[12630], wl[12631], wl[12632], wl[12633], wl[12634], wl[12635], wl[12636], wl[12637], wl[12638], wl[12639], wl[12640], wl[12641], wl[12642], wl[12643], wl[12644], wl[12645], wl[12646], wl[12647], wl[12648], wl[12649], wl[12650], wl[12651], wl[12652], wl[12653], wl[12654], wl[12655], wl[12656], wl[12657], wl[12658], wl[12659], wl[12660], wl[12661], wl[12662], wl[12663], wl[12664], wl[12665], wl[12666], wl[12667], wl[12668], wl[12669], wl[12670], wl[12671], wl[12672], wl[12673], wl[12674], wl[12675], wl[12676], wl[12677], wl[12678], wl[12679], wl[12680], wl[12681], wl[12682], wl[12683], wl[12684], wl[12685], wl[12686], wl[12687], wl[12688], wl[12689], wl[12690], wl[12691], wl[12692], wl[12693], wl[12694], wl[12695], wl[12696], wl[12697], wl[12698], wl[12699], wl[12700], wl[12701], wl[12702], wl[12703], wl[20328], wl[20329], wl[20330], wl[20331], wl[20332], wl[20333], wl[20334], wl[20335], wl[20336], wl[20337], wl[20338], wl[20339], wl[20340], wl[20341], wl[20342], wl[20343], wl[20344], wl[20345], wl[20346], wl[20347], wl[20348], wl[20349], wl[20350], wl[20351], wl[20352], wl[20353], wl[20354], wl[20355], wl[20356], wl[20357], wl[20358], wl[20359], wl[20360], wl[20361], wl[20362], wl[20363], wl[20364], wl[20365], wl[20366], wl[20367], wl[20368], wl[20369], wl[20370], wl[20371], wl[20372], wl[20373], wl[20374], wl[20375], wl[20376], wl[20377], wl[20378], wl[20379], wl[20380], wl[20381], wl[20382], wl[20383], wl[20384], wl[20385], wl[20386], wl[20387], wl[20388], wl[20389], wl[20390], wl[20391], wl[20392], wl[20393], wl[20394], wl[20395], wl[20396], wl[20397], wl[20398], wl[20399], wl[20400], wl[20401], wl[20402], wl[20403], wl[20404], wl[20405], wl[20406], wl[20407], wl[11604], wl[11605], wl[11606], wl[11607], wl[11608], wl[11609], wl[11610], wl[11611], wl[11612], wl[11613], wl[11614], wl[11615], wl[11616], wl[11617], wl[11618], wl[11619], wl[11620], wl[11621], wl[11622], wl[11623], wl[11624], wl[11625], wl[11626], wl[11627], wl[11628], wl[11629], wl[11630], wl[11631], wl[11632], wl[11633], wl[11634], wl[11635], wl[11636], wl[11637], wl[11638], wl[11639], wl[11640], wl[11641], wl[11642], wl[11643], wl[11644], wl[11645], wl[11646], wl[11647], wl[11648], wl[11649], wl[11650], wl[11651], wl[11652], wl[11653], wl[11654], wl[11655], wl[11656], wl[11657], wl[11658], wl[11659], wl[11660], wl[11661], wl[11662], wl[11663], wl[11664], wl[11665], wl[11666], wl[11667], wl[11668], wl[11669], wl[11670], wl[11671], wl[11672], wl[11673], wl[11674], wl[11675], wl[11676], wl[11677], wl[11678], wl[11679], wl[11680], wl[11681], wl[11682], wl[11683], wl[20248], wl[20249], wl[20250], wl[20251], wl[20252], wl[20253], wl[20254], wl[20255], wl[20256], wl[20257], wl[20258], wl[20259], wl[20260], wl[20261], wl[20262], wl[20263], wl[20264], wl[20265], wl[20266], wl[20267], wl[20268], wl[20269], wl[20270], wl[20271], wl[20272], wl[20273], wl[20274], wl[20275], wl[20276], wl[20277], wl[20278], wl[20279], wl[20280], wl[20281], wl[20282], wl[20283], wl[20284], wl[20285], wl[20286], wl[20287], wl[20288], wl[20289], wl[20290], wl[20291], wl[20292], wl[20293], wl[20294], wl[20295], wl[20296], wl[20297], wl[20298], wl[20299], wl[20300], wl[20301], wl[20302], wl[20303], wl[20304], wl[20305], wl[20306], wl[20307], wl[20308], wl[20309], wl[20310], wl[20311], wl[20312], wl[20313], wl[20314], wl[20315], wl[20316], wl[20317], wl[20318], wl[20319], wl[20320], wl[20321], wl[20322], wl[20323], wl[20324], wl[20325], wl[20326], wl[20327]})
    );
    tile tile_3__2_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_1__1__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_1__1__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_1__1__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_2__0__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_2__0__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_2__0__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_1__0__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_1__0__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_1__0__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_1__0__grid_top_r_in[1]),
        .grid_left_in(grid_clb_2__1__grid_left_in),
        .grid_bottom_in(grid_clb_2__1__grid_bottom_in),
        .chanx_left_in(sb_1__1__0_chanx_right_out),
        .chanx_left_out(cbx_1__1__3_chanx_left_out),
        .grid_top_out(grid_clb_2__2__grid_bottom_in),
        .chany_bottom_in(sb_1__0__1_chany_top_out),
        .chany_bottom_out(cby_1__1__4_chany_bottom_out),
        .grid_right_out(grid_clb_3__1__grid_left_in),
        .chany_top_in_0(cby_1__1__5_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__6_chanx_left_out),
        .chany_top_out_0(sb_1__1__3_chany_top_out),
        .chanx_right_out_0(sb_1__1__3_chanx_right_out),
        .grid_top_r_in(sb_2__1__grid_top_r_in),
        .grid_top_l_in(sb_2__1__grid_top_l_in),
        .grid_right_t_in(sb_2__1__grid_right_t_in),
        .grid_right_b_in(sb_2__1__grid_right_b_in),
        .grid_bottom_r_in(sb_2__0__grid_top_r_in),
        .grid_bottom_l_in(sb_2__0__grid_top_l_in),
        .grid_left_t_in(sb_1__1__grid_right_t_in),
        .grid_left_b_in(sb_1__1__grid_right_b_in),
        .bl({bl[2898], bl[2899], bl[2900], bl[2901], bl[2902], bl[2903], bl[2904], bl[2905], bl[2906], bl[2907], bl[2908], bl[2909], bl[2910], bl[2911], bl[2912], bl[2913], bl[2914], bl[2915], bl[2916], bl[2917], bl[2918], bl[2919], bl[2920], bl[2921], bl[2922], bl[2923], bl[2924], bl[2925], bl[2926], bl[2927], bl[2928], bl[2929], bl[2930], bl[2931], bl[2932], bl[2933], bl[2934], bl[2935], bl[2936], bl[2937], bl[2938], bl[2939], bl[2940], bl[2941], bl[2942], bl[2943], bl[2944], bl[2945], bl[2946], bl[2947], bl[2948], bl[2949], bl[2950], bl[2951], bl[2952], bl[2953], bl[2954], bl[2955], bl[2956], bl[2957], bl[2958], bl[2959], bl[2960], bl[2961], bl[2962], bl[2963], bl[2964], bl[2965], bl[2966], bl[2967], bl[2968], bl[2969], bl[2970], bl[2971], bl[2972], bl[2973], bl[2974], bl[2975], bl[2976], bl[2977], bl[2978], bl[2979], bl[2980], bl[2981], bl[2982], bl[2983], bl[2984], bl[2985], bl[2986], bl[2987], bl[2988], bl[2989], bl[2990], bl[2991], bl[2992], bl[2993], bl[2994], bl[2995], bl[2996], bl[2997], bl[2998], bl[2999], bl[3000], bl[3001], bl[3002], bl[3003], bl[3004], bl[3005], bl[3006], bl[3007], bl[3008], bl[3009], bl[3010], bl[3011], bl[3012], bl[3013], bl[3014], bl[3015], bl[3016], bl[3017], bl[3018], bl[3019], bl[3020], bl[3021], bl[3022], bl[3023], bl[3024], bl[3025], bl[3026], bl[3027], bl[3028], bl[3029], bl[3030], bl[3031], bl[3032], bl[3033], bl[3034], bl[3035], bl[3036], bl[3037], bl[3038], bl[3039], bl[3040], bl[3041], bl[3042], bl[3043], bl[3044], bl[3045], bl[3046], bl[3047], bl[3048], bl[3049], bl[3050], bl[3051], bl[3052], bl[3053], bl[3054], bl[3055], bl[3056], bl[3057], bl[3058], bl[3059], bl[3060], bl[3061], bl[3062], bl[3063], bl[3064], bl[3065], bl[3066], bl[3067], bl[3068], bl[3069], bl[3070], bl[3071], bl[3072], bl[3073], bl[3074], bl[3075], bl[3076], bl[3077], bl[3078], bl[3079], bl[3080], bl[3081], bl[3082], bl[3083], bl[3084], bl[3085], bl[3086], bl[3087], bl[3088], bl[3089], bl[3090], bl[3091], bl[3092], bl[3093], bl[3094], bl[3095], bl[3096], bl[3097], bl[3098], bl[3099], bl[3100], bl[3101], bl[3102], bl[3103], bl[3104], bl[3105], bl[3106], bl[3107], bl[3108], bl[3109], bl[3110], bl[3111], bl[3112], bl[3113], bl[3114], bl[3115], bl[3116], bl[3117], bl[3118], bl[3119], bl[3120], bl[3121], bl[3122], bl[3123], bl[3124], bl[3125], bl[3126], bl[3127], bl[3128], bl[3129], bl[3130], bl[3131], bl[3132], bl[3133], bl[3134], bl[3135], bl[3136], bl[3137], bl[3138], bl[3139], bl[3140], bl[3141], bl[3142], bl[3143], bl[3144], bl[3145], bl[3146], bl[3147], bl[3148], bl[3149], bl[3150], bl[3151], bl[3152], bl[3153], bl[3154], bl[3155], bl[3156], bl[3157], bl[3158], bl[3159], bl[3160], bl[3161], bl[3162], bl[3163], bl[3164], bl[3165], bl[3166], bl[3167], bl[3168], bl[3169], bl[3170], bl[3171], bl[3172], bl[3173], bl[3174], bl[3175], bl[3176], bl[3177], bl[3178], bl[3179], bl[3180], bl[3181], bl[3182], bl[3183], bl[3184], bl[3185], bl[3186], bl[3187], bl[3188], bl[3189], bl[3190], bl[3191], bl[3192], bl[3193], bl[3194], bl[3195], bl[3196], bl[3197], bl[3198], bl[3199], bl[3200], bl[3201], bl[3202], bl[3203], bl[3204], bl[3205], bl[3206], bl[3207], bl[3208], bl[3209], bl[3210], bl[3211], bl[3212], bl[3213], bl[3214], bl[3215], bl[3216], bl[3217], bl[3218], bl[3219], bl[3220], bl[3221], bl[3222], bl[3223], bl[3224], bl[3225], bl[3226], bl[3227], bl[3228], bl[3229], bl[3230], bl[3231], bl[3232], bl[3233], bl[3234], bl[3235], bl[3236], bl[3237], bl[3238], bl[3239], bl[3240], bl[3241], bl[3242], bl[3243], bl[3244], bl[3245], bl[3246], bl[3247], bl[3248], bl[3249], bl[3250], bl[3251], bl[3252], bl[3253], bl[3254], bl[3255], bl[3256], bl[3257], bl[3258], bl[3259], bl[3260], bl[3261], bl[3262], bl[3263], bl[3264], bl[3265], bl[3266], bl[3267], bl[3268], bl[3269], bl[3270], bl[3271], bl[3272], bl[3273], bl[3274], bl[3275], bl[3276], bl[3277], bl[3278], bl[3279], bl[3280], bl[3281], bl[3282], bl[3283], bl[3284], bl[3285], bl[3286], bl[3287], bl[3288], bl[3289], bl[3290], bl[3291], bl[3292], bl[3293], bl[3294], bl[3295], bl[3296], bl[3297], bl[3298], bl[3299], bl[3300], bl[3301], bl[3302], bl[3303], bl[3304], bl[3305], bl[3306], bl[3307], bl[3308], bl[3309], bl[3310], bl[3311], bl[3312], bl[3313], bl[3314], bl[3315], bl[3316], bl[3317], bl[3318], bl[3319], bl[3320], bl[3321], bl[3322], bl[3323], bl[3324], bl[3325], bl[3326], bl[3327], bl[3328], bl[3329], bl[3330], bl[3331], bl[3332], bl[3333], bl[3334], bl[3335], bl[3336], bl[3337], bl[3338], bl[3339], bl[3340], bl[3341], bl[3342], bl[3343], bl[3344], bl[3345], bl[3346], bl[3347], bl[3348], bl[3349], bl[3350], bl[3351], bl[3352], bl[3353], bl[3354], bl[3355], bl[3356], bl[3357], bl[3358], bl[3359], bl[3360], bl[3361], bl[3362], bl[3363], bl[3364], bl[3365], bl[3366], bl[3367], bl[3368], bl[3369], bl[3370], bl[3371], bl[3372], bl[3373], bl[3374], bl[3375], bl[3376], bl[3377], bl[3378], bl[3379], bl[3380], bl[3381], bl[3382], bl[3383], bl[3384], bl[3385], bl[3386], bl[3387], bl[3388], bl[3389], bl[3390], bl[3391], bl[3392], bl[3393], bl[3394], bl[3395], bl[3396], bl[3397], bl[3398], bl[3399], bl[3400], bl[3401], bl[3402], bl[3403], bl[3404], bl[3405], bl[3406], bl[3407], bl[3408], bl[3409], bl[3410], bl[3411], bl[3412], bl[3413], bl[3414], bl[3415], bl[3416], bl[3417], bl[3418], bl[3419], bl[3420], bl[3421], bl[3422], bl[3423], bl[3424], bl[3425], bl[3426], bl[3427], bl[3428], bl[3429], bl[3430], bl[3431], bl[3432], bl[3433], bl[3434], bl[3435], bl[3436], bl[3437], bl[3438], bl[3439], bl[3440], bl[3441], bl[3442], bl[3443], bl[3444], bl[3445], bl[3446], bl[3447], bl[3448], bl[3449], bl[3450], bl[3451], bl[3452], bl[3453], bl[3454], bl[3455], bl[3456], bl[3457], bl[3458], bl[3459], bl[3460], bl[3461], bl[3462], bl[3463], bl[3464], bl[3465], bl[3466], bl[3467], bl[3468], bl[3469], bl[3470], bl[3471], bl[3472], bl[3473], bl[3474], bl[3475], bl[3476], bl[3477], bl[3478], bl[3479], bl[3480], bl[3481], bl[3482], bl[3483], bl[3484], bl[3485], bl[3486], bl[3487], bl[3488], bl[3489], bl[3490], bl[3491], bl[3492], bl[3493], bl[3494], bl[3495], bl[3496], bl[3497], bl[3498], bl[3499], bl[3500], bl[3501], bl[3502], bl[3503], bl[3504], bl[3505], bl[3506], bl[3507], bl[3508], bl[3509], bl[3510], bl[3511], bl[3512], bl[3513], bl[3514], bl[3515], bl[3516], bl[3517], bl[3518], bl[3519], bl[3520], bl[3521], bl[3522], bl[3523], bl[3524], bl[3525], bl[3526], bl[3527], bl[3528], bl[3529], bl[3530], bl[3531], bl[3532], bl[3533], bl[3534], bl[3535], bl[3536], bl[3537], bl[3538], bl[3539], bl[3540], bl[3541], bl[3542], bl[3543], bl[3544], bl[3545], bl[3546], bl[3547], bl[3548], bl[3549], bl[3550], bl[3551], bl[3552], bl[3553], bl[3554], bl[3555], bl[3556], bl[3557], bl[3558], bl[3559], bl[3560], bl[3561], bl[3562], bl[3563], bl[3564], bl[3565], bl[3566], bl[3567], bl[3568], bl[3569], bl[3570], bl[3571], bl[3572], bl[3573], bl[3574], bl[3575], bl[3576], bl[3577], bl[3578], bl[3579], bl[3580], bl[3581], bl[3582], bl[3583], bl[3584], bl[3585], bl[3586], bl[3587], bl[3588], bl[3589], bl[3590], bl[3591], bl[3592], bl[3593], bl[3594], bl[3595], bl[3596], bl[3597], bl[3598], bl[3599], bl[3600], bl[3601], bl[3602], bl[3603], bl[3604], bl[3605], bl[3606], bl[3607], bl[3608], bl[3609], bl[3610], bl[3611], bl[3612], bl[3613], bl[3614], bl[3615], bl[3616], bl[3617], bl[3618], bl[3619], bl[3620], bl[3621], bl[3622], bl[3623], bl[3624], bl[3625], bl[3626], bl[3627], bl[3628], bl[3629], bl[3630], bl[3631], bl[3632], bl[3633], bl[3634], bl[3635], bl[3636], bl[3637], bl[3638], bl[3639], bl[3640], bl[3641], bl[3642], bl[3643], bl[3644], bl[3645], bl[3646], bl[3647], bl[3648], bl[3649], bl[3650], bl[3651], bl[3652], bl[3653], bl[3654], bl[3655], bl[3656], bl[3657], bl[3658], bl[3659], bl[3660], bl[3661], bl[3662], bl[3663], bl[3664], bl[3665], bl[3666], bl[3667], bl[3668], bl[3669], bl[3670], bl[3671], bl[3672], bl[3673], bl[3674], bl[3675], bl[3676], bl[3677], bl[3678], bl[3679], bl[3680], bl[3681], bl[3682], bl[3683], bl[3684], bl[3685], bl[3686], bl[3687], bl[3688], bl[3689], bl[3690], bl[3691], bl[3692], bl[3693], bl[3694], bl[3695], bl[3696], bl[3697], bl[3698], bl[3699], bl[3700], bl[3701], bl[3702], bl[3703], bl[3704], bl[3705], bl[3706], bl[3707], bl[3708], bl[3709], bl[3710], bl[3711], bl[3712], bl[3713], bl[3714], bl[3715], bl[3716], bl[3717], bl[3718], bl[3719], bl[3720], bl[3721], bl[3722], bl[3723], bl[3724], bl[3725], bl[3726], bl[3727], bl[3728], bl[3729], bl[3730], bl[3731], bl[3732], bl[3733], bl[3734], bl[3735], bl[3736], bl[3737], bl[3738], bl[3739], bl[3740], bl[3741], bl[3742], bl[3743], bl[3744], bl[3745], bl[3746], bl[3747], bl[3748], bl[3749], bl[3750], bl[3751], bl[3752], bl[3753], bl[3754], bl[3755], bl[3756], bl[3757], bl[3758], bl[3759], bl[3760], bl[3761], bl[3762], bl[3763], bl[3764], bl[3765], bl[3766], bl[3767], bl[3768], bl[3769], bl[3770], bl[3771], bl[3772], bl[3773], bl[3774], bl[3775], bl[3776], bl[3777], bl[3778], bl[3779], bl[3780], bl[3781], bl[3782], bl[3783], bl[3784], bl[3785], bl[3786], bl[3787], bl[3788], bl[3789], bl[3790], bl[3791], bl[3792], bl[3793], bl[3794], bl[3795], bl[3796], bl[3797], bl[3798], bl[3799], bl[3800], bl[3801], bl[3802], bl[3803], bl[3804], bl[3805], bl[3806], bl[3807], bl[3808], bl[3809], bl[3810], bl[3811], bl[3812], bl[3813], bl[3814], bl[3815], bl[3816], bl[3817], bl[3818], bl[3819], bl[3820], bl[3821], bl[3822], bl[3823], bl[3824], bl[3825], bl[3826], bl[3827], bl[3828], bl[3829], bl[3830], bl[3831], bl[3832], bl[3833], bl[3834], bl[3835], bl[3836], bl[3837], bl[3838], bl[3839], bl[3840], bl[3841], bl[3842], bl[3843], bl[3844], bl[3845], bl[3846], bl[3847], bl[3848], bl[3849], bl[3850], bl[3851], bl[3852], bl[3853], bl[3854], bl[3855], bl[3856], bl[3857], bl[3858], bl[3859], bl[3860], bl[3861], bl[3862], bl[3863], bl[3864], bl[3865], bl[3866], bl[3867], bl[3868], bl[3869], bl[3870], bl[3871], bl[3872], bl[3873], bl[3874], bl[3875], bl[3876], bl[3877], bl[3878], bl[3879], bl[3880], bl[3881], bl[3882], bl[3883], bl[3884], bl[3885], bl[3886], bl[3887], bl[3888], bl[3889], bl[3890], bl[3891], bl[3892], bl[3893], bl[3894], bl[3895], bl[3896], bl[3897], bl[3898], bl[3899], bl[3900], bl[3901], bl[3902], bl[3903], bl[3904], bl[3905], bl[3906], bl[3907], bl[3908], bl[3909], bl[3910], bl[3911], bl[3912], bl[3913], bl[3914], bl[3915], bl[3916], bl[3917], bl[9004], bl[9005], bl[9006], bl[9007], bl[9008], bl[9009], bl[9010], bl[9011], bl[9012], bl[9013], bl[9014], bl[9015], bl[9016], bl[9017], bl[9018], bl[9019], bl[9020], bl[9021], bl[9022], bl[9023], bl[9024], bl[9025], bl[9026], bl[9027], bl[9028], bl[9029], bl[9030], bl[9031], bl[9032], bl[9033], bl[9034], bl[9035], bl[9036], bl[9037], bl[9038], bl[9039], bl[9040], bl[9041], bl[9042], bl[9043], bl[9044], bl[9045], bl[9046], bl[9047], bl[9048], bl[9049], bl[9050], bl[9051], bl[9052], bl[9053], bl[9054], bl[9055], bl[9056], bl[9057], bl[9058], bl[9059], bl[9060], bl[9061], bl[9062], bl[9063], bl[9064], bl[9065], bl[9066], bl[9067], bl[9068], bl[9069], bl[9070], bl[9071], bl[9072], bl[9073], bl[9074], bl[9075], bl[9076], bl[9077], bl[9078], bl[9079], bl[9080], bl[9081], bl[9082], bl[9083], bl[2818], bl[2819], bl[2820], bl[2821], bl[2822], bl[2823], bl[2824], bl[2825], bl[2826], bl[2827], bl[2828], bl[2829], bl[2830], bl[2831], bl[2832], bl[2833], bl[2834], bl[2835], bl[2836], bl[2837], bl[2838], bl[2839], bl[2840], bl[2841], bl[2842], bl[2843], bl[2844], bl[2845], bl[2846], bl[2847], bl[2848], bl[2849], bl[2850], bl[2851], bl[2852], bl[2853], bl[2854], bl[2855], bl[2856], bl[2857], bl[2858], bl[2859], bl[2860], bl[2861], bl[2862], bl[2863], bl[2864], bl[2865], bl[2866], bl[2867], bl[2868], bl[2869], bl[2870], bl[2871], bl[2872], bl[2873], bl[2874], bl[2875], bl[2876], bl[2877], bl[2878], bl[2879], bl[2880], bl[2881], bl[2882], bl[2883], bl[2884], bl[2885], bl[2886], bl[2887], bl[2888], bl[2889], bl[2890], bl[2891], bl[2892], bl[2893], bl[2894], bl[2895], bl[2896], bl[2897], bl[8924], bl[8925], bl[8926], bl[8927], bl[8928], bl[8929], bl[8930], bl[8931], bl[8932], bl[8933], bl[8934], bl[8935], bl[8936], bl[8937], bl[8938], bl[8939], bl[8940], bl[8941], bl[8942], bl[8943], bl[8944], bl[8945], bl[8946], bl[8947], bl[8948], bl[8949], bl[8950], bl[8951], bl[8952], bl[8953], bl[8954], bl[8955], bl[8956], bl[8957], bl[8958], bl[8959], bl[8960], bl[8961], bl[8962], bl[8963], bl[8964], bl[8965], bl[8966], bl[8967], bl[8968], bl[8969], bl[8970], bl[8971], bl[8972], bl[8973], bl[8974], bl[8975], bl[8976], bl[8977], bl[8978], bl[8979], bl[8980], bl[8981], bl[8982], bl[8983], bl[8984], bl[8985], bl[8986], bl[8987], bl[8988], bl[8989], bl[8990], bl[8991], bl[8992], bl[8993], bl[8994], bl[8995], bl[8996], bl[8997], bl[8998], bl[8999], bl[9000], bl[9001], bl[9002], bl[9003]}),
        .wl({wl[2898], wl[2899], wl[2900], wl[2901], wl[2902], wl[2903], wl[2904], wl[2905], wl[2906], wl[2907], wl[2908], wl[2909], wl[2910], wl[2911], wl[2912], wl[2913], wl[2914], wl[2915], wl[2916], wl[2917], wl[2918], wl[2919], wl[2920], wl[2921], wl[2922], wl[2923], wl[2924], wl[2925], wl[2926], wl[2927], wl[2928], wl[2929], wl[2930], wl[2931], wl[2932], wl[2933], wl[2934], wl[2935], wl[2936], wl[2937], wl[2938], wl[2939], wl[2940], wl[2941], wl[2942], wl[2943], wl[2944], wl[2945], wl[2946], wl[2947], wl[2948], wl[2949], wl[2950], wl[2951], wl[2952], wl[2953], wl[2954], wl[2955], wl[2956], wl[2957], wl[2958], wl[2959], wl[2960], wl[2961], wl[2962], wl[2963], wl[2964], wl[2965], wl[2966], wl[2967], wl[2968], wl[2969], wl[2970], wl[2971], wl[2972], wl[2973], wl[2974], wl[2975], wl[2976], wl[2977], wl[2978], wl[2979], wl[2980], wl[2981], wl[2982], wl[2983], wl[2984], wl[2985], wl[2986], wl[2987], wl[2988], wl[2989], wl[2990], wl[2991], wl[2992], wl[2993], wl[2994], wl[2995], wl[2996], wl[2997], wl[2998], wl[2999], wl[3000], wl[3001], wl[3002], wl[3003], wl[3004], wl[3005], wl[3006], wl[3007], wl[3008], wl[3009], wl[3010], wl[3011], wl[3012], wl[3013], wl[3014], wl[3015], wl[3016], wl[3017], wl[3018], wl[3019], wl[3020], wl[3021], wl[3022], wl[3023], wl[3024], wl[3025], wl[3026], wl[3027], wl[3028], wl[3029], wl[3030], wl[3031], wl[3032], wl[3033], wl[3034], wl[3035], wl[3036], wl[3037], wl[3038], wl[3039], wl[3040], wl[3041], wl[3042], wl[3043], wl[3044], wl[3045], wl[3046], wl[3047], wl[3048], wl[3049], wl[3050], wl[3051], wl[3052], wl[3053], wl[3054], wl[3055], wl[3056], wl[3057], wl[3058], wl[3059], wl[3060], wl[3061], wl[3062], wl[3063], wl[3064], wl[3065], wl[3066], wl[3067], wl[3068], wl[3069], wl[3070], wl[3071], wl[3072], wl[3073], wl[3074], wl[3075], wl[3076], wl[3077], wl[3078], wl[3079], wl[3080], wl[3081], wl[3082], wl[3083], wl[3084], wl[3085], wl[3086], wl[3087], wl[3088], wl[3089], wl[3090], wl[3091], wl[3092], wl[3093], wl[3094], wl[3095], wl[3096], wl[3097], wl[3098], wl[3099], wl[3100], wl[3101], wl[3102], wl[3103], wl[3104], wl[3105], wl[3106], wl[3107], wl[3108], wl[3109], wl[3110], wl[3111], wl[3112], wl[3113], wl[3114], wl[3115], wl[3116], wl[3117], wl[3118], wl[3119], wl[3120], wl[3121], wl[3122], wl[3123], wl[3124], wl[3125], wl[3126], wl[3127], wl[3128], wl[3129], wl[3130], wl[3131], wl[3132], wl[3133], wl[3134], wl[3135], wl[3136], wl[3137], wl[3138], wl[3139], wl[3140], wl[3141], wl[3142], wl[3143], wl[3144], wl[3145], wl[3146], wl[3147], wl[3148], wl[3149], wl[3150], wl[3151], wl[3152], wl[3153], wl[3154], wl[3155], wl[3156], wl[3157], wl[3158], wl[3159], wl[3160], wl[3161], wl[3162], wl[3163], wl[3164], wl[3165], wl[3166], wl[3167], wl[3168], wl[3169], wl[3170], wl[3171], wl[3172], wl[3173], wl[3174], wl[3175], wl[3176], wl[3177], wl[3178], wl[3179], wl[3180], wl[3181], wl[3182], wl[3183], wl[3184], wl[3185], wl[3186], wl[3187], wl[3188], wl[3189], wl[3190], wl[3191], wl[3192], wl[3193], wl[3194], wl[3195], wl[3196], wl[3197], wl[3198], wl[3199], wl[3200], wl[3201], wl[3202], wl[3203], wl[3204], wl[3205], wl[3206], wl[3207], wl[3208], wl[3209], wl[3210], wl[3211], wl[3212], wl[3213], wl[3214], wl[3215], wl[3216], wl[3217], wl[3218], wl[3219], wl[3220], wl[3221], wl[3222], wl[3223], wl[3224], wl[3225], wl[3226], wl[3227], wl[3228], wl[3229], wl[3230], wl[3231], wl[3232], wl[3233], wl[3234], wl[3235], wl[3236], wl[3237], wl[3238], wl[3239], wl[3240], wl[3241], wl[3242], wl[3243], wl[3244], wl[3245], wl[3246], wl[3247], wl[3248], wl[3249], wl[3250], wl[3251], wl[3252], wl[3253], wl[3254], wl[3255], wl[3256], wl[3257], wl[3258], wl[3259], wl[3260], wl[3261], wl[3262], wl[3263], wl[3264], wl[3265], wl[3266], wl[3267], wl[3268], wl[3269], wl[3270], wl[3271], wl[3272], wl[3273], wl[3274], wl[3275], wl[3276], wl[3277], wl[3278], wl[3279], wl[3280], wl[3281], wl[3282], wl[3283], wl[3284], wl[3285], wl[3286], wl[3287], wl[3288], wl[3289], wl[3290], wl[3291], wl[3292], wl[3293], wl[3294], wl[3295], wl[3296], wl[3297], wl[3298], wl[3299], wl[3300], wl[3301], wl[3302], wl[3303], wl[3304], wl[3305], wl[3306], wl[3307], wl[3308], wl[3309], wl[3310], wl[3311], wl[3312], wl[3313], wl[3314], wl[3315], wl[3316], wl[3317], wl[3318], wl[3319], wl[3320], wl[3321], wl[3322], wl[3323], wl[3324], wl[3325], wl[3326], wl[3327], wl[3328], wl[3329], wl[3330], wl[3331], wl[3332], wl[3333], wl[3334], wl[3335], wl[3336], wl[3337], wl[3338], wl[3339], wl[3340], wl[3341], wl[3342], wl[3343], wl[3344], wl[3345], wl[3346], wl[3347], wl[3348], wl[3349], wl[3350], wl[3351], wl[3352], wl[3353], wl[3354], wl[3355], wl[3356], wl[3357], wl[3358], wl[3359], wl[3360], wl[3361], wl[3362], wl[3363], wl[3364], wl[3365], wl[3366], wl[3367], wl[3368], wl[3369], wl[3370], wl[3371], wl[3372], wl[3373], wl[3374], wl[3375], wl[3376], wl[3377], wl[3378], wl[3379], wl[3380], wl[3381], wl[3382], wl[3383], wl[3384], wl[3385], wl[3386], wl[3387], wl[3388], wl[3389], wl[3390], wl[3391], wl[3392], wl[3393], wl[3394], wl[3395], wl[3396], wl[3397], wl[3398], wl[3399], wl[3400], wl[3401], wl[3402], wl[3403], wl[3404], wl[3405], wl[3406], wl[3407], wl[3408], wl[3409], wl[3410], wl[3411], wl[3412], wl[3413], wl[3414], wl[3415], wl[3416], wl[3417], wl[3418], wl[3419], wl[3420], wl[3421], wl[3422], wl[3423], wl[3424], wl[3425], wl[3426], wl[3427], wl[3428], wl[3429], wl[3430], wl[3431], wl[3432], wl[3433], wl[3434], wl[3435], wl[3436], wl[3437], wl[3438], wl[3439], wl[3440], wl[3441], wl[3442], wl[3443], wl[3444], wl[3445], wl[3446], wl[3447], wl[3448], wl[3449], wl[3450], wl[3451], wl[3452], wl[3453], wl[3454], wl[3455], wl[3456], wl[3457], wl[3458], wl[3459], wl[3460], wl[3461], wl[3462], wl[3463], wl[3464], wl[3465], wl[3466], wl[3467], wl[3468], wl[3469], wl[3470], wl[3471], wl[3472], wl[3473], wl[3474], wl[3475], wl[3476], wl[3477], wl[3478], wl[3479], wl[3480], wl[3481], wl[3482], wl[3483], wl[3484], wl[3485], wl[3486], wl[3487], wl[3488], wl[3489], wl[3490], wl[3491], wl[3492], wl[3493], wl[3494], wl[3495], wl[3496], wl[3497], wl[3498], wl[3499], wl[3500], wl[3501], wl[3502], wl[3503], wl[3504], wl[3505], wl[3506], wl[3507], wl[3508], wl[3509], wl[3510], wl[3511], wl[3512], wl[3513], wl[3514], wl[3515], wl[3516], wl[3517], wl[3518], wl[3519], wl[3520], wl[3521], wl[3522], wl[3523], wl[3524], wl[3525], wl[3526], wl[3527], wl[3528], wl[3529], wl[3530], wl[3531], wl[3532], wl[3533], wl[3534], wl[3535], wl[3536], wl[3537], wl[3538], wl[3539], wl[3540], wl[3541], wl[3542], wl[3543], wl[3544], wl[3545], wl[3546], wl[3547], wl[3548], wl[3549], wl[3550], wl[3551], wl[3552], wl[3553], wl[3554], wl[3555], wl[3556], wl[3557], wl[3558], wl[3559], wl[3560], wl[3561], wl[3562], wl[3563], wl[3564], wl[3565], wl[3566], wl[3567], wl[3568], wl[3569], wl[3570], wl[3571], wl[3572], wl[3573], wl[3574], wl[3575], wl[3576], wl[3577], wl[3578], wl[3579], wl[3580], wl[3581], wl[3582], wl[3583], wl[3584], wl[3585], wl[3586], wl[3587], wl[3588], wl[3589], wl[3590], wl[3591], wl[3592], wl[3593], wl[3594], wl[3595], wl[3596], wl[3597], wl[3598], wl[3599], wl[3600], wl[3601], wl[3602], wl[3603], wl[3604], wl[3605], wl[3606], wl[3607], wl[3608], wl[3609], wl[3610], wl[3611], wl[3612], wl[3613], wl[3614], wl[3615], wl[3616], wl[3617], wl[3618], wl[3619], wl[3620], wl[3621], wl[3622], wl[3623], wl[3624], wl[3625], wl[3626], wl[3627], wl[3628], wl[3629], wl[3630], wl[3631], wl[3632], wl[3633], wl[3634], wl[3635], wl[3636], wl[3637], wl[3638], wl[3639], wl[3640], wl[3641], wl[3642], wl[3643], wl[3644], wl[3645], wl[3646], wl[3647], wl[3648], wl[3649], wl[3650], wl[3651], wl[3652], wl[3653], wl[3654], wl[3655], wl[3656], wl[3657], wl[3658], wl[3659], wl[3660], wl[3661], wl[3662], wl[3663], wl[3664], wl[3665], wl[3666], wl[3667], wl[3668], wl[3669], wl[3670], wl[3671], wl[3672], wl[3673], wl[3674], wl[3675], wl[3676], wl[3677], wl[3678], wl[3679], wl[3680], wl[3681], wl[3682], wl[3683], wl[3684], wl[3685], wl[3686], wl[3687], wl[3688], wl[3689], wl[3690], wl[3691], wl[3692], wl[3693], wl[3694], wl[3695], wl[3696], wl[3697], wl[3698], wl[3699], wl[3700], wl[3701], wl[3702], wl[3703], wl[3704], wl[3705], wl[3706], wl[3707], wl[3708], wl[3709], wl[3710], wl[3711], wl[3712], wl[3713], wl[3714], wl[3715], wl[3716], wl[3717], wl[3718], wl[3719], wl[3720], wl[3721], wl[3722], wl[3723], wl[3724], wl[3725], wl[3726], wl[3727], wl[3728], wl[3729], wl[3730], wl[3731], wl[3732], wl[3733], wl[3734], wl[3735], wl[3736], wl[3737], wl[3738], wl[3739], wl[3740], wl[3741], wl[3742], wl[3743], wl[3744], wl[3745], wl[3746], wl[3747], wl[3748], wl[3749], wl[3750], wl[3751], wl[3752], wl[3753], wl[3754], wl[3755], wl[3756], wl[3757], wl[3758], wl[3759], wl[3760], wl[3761], wl[3762], wl[3763], wl[3764], wl[3765], wl[3766], wl[3767], wl[3768], wl[3769], wl[3770], wl[3771], wl[3772], wl[3773], wl[3774], wl[3775], wl[3776], wl[3777], wl[3778], wl[3779], wl[3780], wl[3781], wl[3782], wl[3783], wl[3784], wl[3785], wl[3786], wl[3787], wl[3788], wl[3789], wl[3790], wl[3791], wl[3792], wl[3793], wl[3794], wl[3795], wl[3796], wl[3797], wl[3798], wl[3799], wl[3800], wl[3801], wl[3802], wl[3803], wl[3804], wl[3805], wl[3806], wl[3807], wl[3808], wl[3809], wl[3810], wl[3811], wl[3812], wl[3813], wl[3814], wl[3815], wl[3816], wl[3817], wl[3818], wl[3819], wl[3820], wl[3821], wl[3822], wl[3823], wl[3824], wl[3825], wl[3826], wl[3827], wl[3828], wl[3829], wl[3830], wl[3831], wl[3832], wl[3833], wl[3834], wl[3835], wl[3836], wl[3837], wl[3838], wl[3839], wl[3840], wl[3841], wl[3842], wl[3843], wl[3844], wl[3845], wl[3846], wl[3847], wl[3848], wl[3849], wl[3850], wl[3851], wl[3852], wl[3853], wl[3854], wl[3855], wl[3856], wl[3857], wl[3858], wl[3859], wl[3860], wl[3861], wl[3862], wl[3863], wl[3864], wl[3865], wl[3866], wl[3867], wl[3868], wl[3869], wl[3870], wl[3871], wl[3872], wl[3873], wl[3874], wl[3875], wl[3876], wl[3877], wl[3878], wl[3879], wl[3880], wl[3881], wl[3882], wl[3883], wl[3884], wl[3885], wl[3886], wl[3887], wl[3888], wl[3889], wl[3890], wl[3891], wl[3892], wl[3893], wl[3894], wl[3895], wl[3896], wl[3897], wl[3898], wl[3899], wl[3900], wl[3901], wl[3902], wl[3903], wl[3904], wl[3905], wl[3906], wl[3907], wl[3908], wl[3909], wl[3910], wl[3911], wl[3912], wl[3913], wl[3914], wl[3915], wl[3916], wl[3917], wl[9004], wl[9005], wl[9006], wl[9007], wl[9008], wl[9009], wl[9010], wl[9011], wl[9012], wl[9013], wl[9014], wl[9015], wl[9016], wl[9017], wl[9018], wl[9019], wl[9020], wl[9021], wl[9022], wl[9023], wl[9024], wl[9025], wl[9026], wl[9027], wl[9028], wl[9029], wl[9030], wl[9031], wl[9032], wl[9033], wl[9034], wl[9035], wl[9036], wl[9037], wl[9038], wl[9039], wl[9040], wl[9041], wl[9042], wl[9043], wl[9044], wl[9045], wl[9046], wl[9047], wl[9048], wl[9049], wl[9050], wl[9051], wl[9052], wl[9053], wl[9054], wl[9055], wl[9056], wl[9057], wl[9058], wl[9059], wl[9060], wl[9061], wl[9062], wl[9063], wl[9064], wl[9065], wl[9066], wl[9067], wl[9068], wl[9069], wl[9070], wl[9071], wl[9072], wl[9073], wl[9074], wl[9075], wl[9076], wl[9077], wl[9078], wl[9079], wl[9080], wl[9081], wl[9082], wl[9083], wl[2818], wl[2819], wl[2820], wl[2821], wl[2822], wl[2823], wl[2824], wl[2825], wl[2826], wl[2827], wl[2828], wl[2829], wl[2830], wl[2831], wl[2832], wl[2833], wl[2834], wl[2835], wl[2836], wl[2837], wl[2838], wl[2839], wl[2840], wl[2841], wl[2842], wl[2843], wl[2844], wl[2845], wl[2846], wl[2847], wl[2848], wl[2849], wl[2850], wl[2851], wl[2852], wl[2853], wl[2854], wl[2855], wl[2856], wl[2857], wl[2858], wl[2859], wl[2860], wl[2861], wl[2862], wl[2863], wl[2864], wl[2865], wl[2866], wl[2867], wl[2868], wl[2869], wl[2870], wl[2871], wl[2872], wl[2873], wl[2874], wl[2875], wl[2876], wl[2877], wl[2878], wl[2879], wl[2880], wl[2881], wl[2882], wl[2883], wl[2884], wl[2885], wl[2886], wl[2887], wl[2888], wl[2889], wl[2890], wl[2891], wl[2892], wl[2893], wl[2894], wl[2895], wl[2896], wl[2897], wl[8924], wl[8925], wl[8926], wl[8927], wl[8928], wl[8929], wl[8930], wl[8931], wl[8932], wl[8933], wl[8934], wl[8935], wl[8936], wl[8937], wl[8938], wl[8939], wl[8940], wl[8941], wl[8942], wl[8943], wl[8944], wl[8945], wl[8946], wl[8947], wl[8948], wl[8949], wl[8950], wl[8951], wl[8952], wl[8953], wl[8954], wl[8955], wl[8956], wl[8957], wl[8958], wl[8959], wl[8960], wl[8961], wl[8962], wl[8963], wl[8964], wl[8965], wl[8966], wl[8967], wl[8968], wl[8969], wl[8970], wl[8971], wl[8972], wl[8973], wl[8974], wl[8975], wl[8976], wl[8977], wl[8978], wl[8979], wl[8980], wl[8981], wl[8982], wl[8983], wl[8984], wl[8985], wl[8986], wl[8987], wl[8988], wl[8989], wl[8990], wl[8991], wl[8992], wl[8993], wl[8994], wl[8995], wl[8996], wl[8997], wl[8998], wl[8999], wl[9000], wl[9001], wl[9002], wl[9003]})
    );
    tile tile_3__3_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_1__2__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_1__2__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_1__2__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_2__1__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_2__1__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_2__1__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_1__1__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_1__1__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_1__1__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_1__1__grid_top_r_in[1]),
        .grid_left_in(grid_clb_2__2__grid_left_in),
        .grid_bottom_in(grid_clb_2__2__grid_bottom_in),
        .chanx_left_in(sb_1__1__1_chanx_right_out),
        .chanx_left_out(cbx_1__1__4_chanx_left_out),
        .grid_top_out(grid_clb_2__3__grid_bottom_in),
        .chany_bottom_in(sb_1__1__3_chany_top_out),
        .chany_bottom_out(cby_1__1__5_chany_bottom_out),
        .grid_right_out(grid_clb_3__2__grid_left_in),
        .chany_top_in_0(cby_1__1__6_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__7_chanx_left_out),
        .chany_top_out_0(sb_1__1__4_chany_top_out),
        .chanx_right_out_0(sb_1__1__4_chanx_right_out),
        .grid_top_r_in(sb_2__2__grid_top_r_in),
        .grid_top_l_in(sb_2__2__grid_top_l_in),
        .grid_right_t_in(sb_2__2__grid_right_t_in),
        .grid_right_b_in(sb_2__2__grid_right_b_in),
        .grid_bottom_r_in(sb_2__1__grid_top_r_in),
        .grid_bottom_l_in(sb_2__1__grid_top_l_in),
        .grid_left_t_in(sb_1__2__grid_right_t_in),
        .grid_left_b_in(sb_1__2__grid_right_b_in),
        .bl({bl[9164], bl[9165], bl[9166], bl[9167], bl[9168], bl[9169], bl[9170], bl[9171], bl[9172], bl[9173], bl[9174], bl[9175], bl[9176], bl[9177], bl[9178], bl[9179], bl[9180], bl[9181], bl[9182], bl[9183], bl[9184], bl[9185], bl[9186], bl[9187], bl[9188], bl[9189], bl[9190], bl[9191], bl[9192], bl[9193], bl[9194], bl[9195], bl[9196], bl[9197], bl[9198], bl[9199], bl[9200], bl[9201], bl[9202], bl[9203], bl[9204], bl[9205], bl[9206], bl[9207], bl[9208], bl[9209], bl[9210], bl[9211], bl[9212], bl[9213], bl[9214], bl[9215], bl[9216], bl[9217], bl[9218], bl[9219], bl[9220], bl[9221], bl[9222], bl[9223], bl[9224], bl[9225], bl[9226], bl[9227], bl[9228], bl[9229], bl[9230], bl[9231], bl[9232], bl[9233], bl[9234], bl[9235], bl[9236], bl[9237], bl[9238], bl[9239], bl[9240], bl[9241], bl[9242], bl[9243], bl[9244], bl[9245], bl[9246], bl[9247], bl[9248], bl[9249], bl[9250], bl[9251], bl[9252], bl[9253], bl[9254], bl[9255], bl[9256], bl[9257], bl[9258], bl[9259], bl[9260], bl[9261], bl[9262], bl[9263], bl[9264], bl[9265], bl[9266], bl[9267], bl[9268], bl[9269], bl[9270], bl[9271], bl[9272], bl[9273], bl[9274], bl[9275], bl[9276], bl[9277], bl[9278], bl[9279], bl[9280], bl[9281], bl[9282], bl[9283], bl[9284], bl[9285], bl[9286], bl[9287], bl[9288], bl[9289], bl[9290], bl[9291], bl[9292], bl[9293], bl[9294], bl[9295], bl[9296], bl[9297], bl[9298], bl[9299], bl[9300], bl[9301], bl[9302], bl[9303], bl[9304], bl[9305], bl[9306], bl[9307], bl[9308], bl[9309], bl[9310], bl[9311], bl[9312], bl[9313], bl[9314], bl[9315], bl[9316], bl[9317], bl[9318], bl[9319], bl[9320], bl[9321], bl[9322], bl[9323], bl[9324], bl[9325], bl[9326], bl[9327], bl[9328], bl[9329], bl[9330], bl[9331], bl[9332], bl[9333], bl[9334], bl[9335], bl[9336], bl[9337], bl[9338], bl[9339], bl[9340], bl[9341], bl[9342], bl[9343], bl[9344], bl[9345], bl[9346], bl[9347], bl[9348], bl[9349], bl[9350], bl[9351], bl[9352], bl[9353], bl[9354], bl[9355], bl[9356], bl[9357], bl[9358], bl[9359], bl[9360], bl[9361], bl[9362], bl[9363], bl[9364], bl[9365], bl[9366], bl[9367], bl[9368], bl[9369], bl[9370], bl[9371], bl[9372], bl[9373], bl[9374], bl[9375], bl[9376], bl[9377], bl[9378], bl[9379], bl[9380], bl[9381], bl[9382], bl[9383], bl[9384], bl[9385], bl[9386], bl[9387], bl[9388], bl[9389], bl[9390], bl[9391], bl[9392], bl[9393], bl[9394], bl[9395], bl[9396], bl[9397], bl[9398], bl[9399], bl[9400], bl[9401], bl[9402], bl[9403], bl[9404], bl[9405], bl[9406], bl[9407], bl[9408], bl[9409], bl[9410], bl[9411], bl[9412], bl[9413], bl[9414], bl[9415], bl[9416], bl[9417], bl[9418], bl[9419], bl[9420], bl[9421], bl[9422], bl[9423], bl[9424], bl[9425], bl[9426], bl[9427], bl[9428], bl[9429], bl[9430], bl[9431], bl[9432], bl[9433], bl[9434], bl[9435], bl[9436], bl[9437], bl[9438], bl[9439], bl[9440], bl[9441], bl[9442], bl[9443], bl[9444], bl[9445], bl[9446], bl[9447], bl[9448], bl[9449], bl[9450], bl[9451], bl[9452], bl[9453], bl[9454], bl[9455], bl[9456], bl[9457], bl[9458], bl[9459], bl[9460], bl[9461], bl[9462], bl[9463], bl[9464], bl[9465], bl[9466], bl[9467], bl[9468], bl[9469], bl[9470], bl[9471], bl[9472], bl[9473], bl[9474], bl[9475], bl[9476], bl[9477], bl[9478], bl[9479], bl[9480], bl[9481], bl[9482], bl[9483], bl[9484], bl[9485], bl[9486], bl[9487], bl[9488], bl[9489], bl[9490], bl[9491], bl[9492], bl[9493], bl[9494], bl[9495], bl[9496], bl[9497], bl[9498], bl[9499], bl[9500], bl[9501], bl[9502], bl[9503], bl[9504], bl[9505], bl[9506], bl[9507], bl[9508], bl[9509], bl[9510], bl[9511], bl[9512], bl[9513], bl[9514], bl[9515], bl[9516], bl[9517], bl[9518], bl[9519], bl[9520], bl[9521], bl[9522], bl[9523], bl[9524], bl[9525], bl[9526], bl[9527], bl[9528], bl[9529], bl[9530], bl[9531], bl[9532], bl[9533], bl[9534], bl[9535], bl[9536], bl[9537], bl[9538], bl[9539], bl[9540], bl[9541], bl[9542], bl[9543], bl[9544], bl[9545], bl[9546], bl[9547], bl[9548], bl[9549], bl[9550], bl[9551], bl[9552], bl[9553], bl[9554], bl[9555], bl[9556], bl[9557], bl[9558], bl[9559], bl[9560], bl[9561], bl[9562], bl[9563], bl[9564], bl[9565], bl[9566], bl[9567], bl[9568], bl[9569], bl[9570], bl[9571], bl[9572], bl[9573], bl[9574], bl[9575], bl[9576], bl[9577], bl[9578], bl[9579], bl[9580], bl[9581], bl[9582], bl[9583], bl[9584], bl[9585], bl[9586], bl[9587], bl[9588], bl[9589], bl[9590], bl[9591], bl[9592], bl[9593], bl[9594], bl[9595], bl[9596], bl[9597], bl[9598], bl[9599], bl[9600], bl[9601], bl[9602], bl[9603], bl[9604], bl[9605], bl[9606], bl[9607], bl[9608], bl[9609], bl[9610], bl[9611], bl[9612], bl[9613], bl[9614], bl[9615], bl[9616], bl[9617], bl[9618], bl[9619], bl[9620], bl[9621], bl[9622], bl[9623], bl[9624], bl[9625], bl[9626], bl[9627], bl[9628], bl[9629], bl[9630], bl[9631], bl[9632], bl[9633], bl[9634], bl[9635], bl[9636], bl[9637], bl[9638], bl[9639], bl[9640], bl[9641], bl[9642], bl[9643], bl[9644], bl[9645], bl[9646], bl[9647], bl[9648], bl[9649], bl[9650], bl[9651], bl[9652], bl[9653], bl[9654], bl[9655], bl[9656], bl[9657], bl[9658], bl[9659], bl[9660], bl[9661], bl[9662], bl[9663], bl[9664], bl[9665], bl[9666], bl[9667], bl[9668], bl[9669], bl[9670], bl[9671], bl[9672], bl[9673], bl[9674], bl[9675], bl[9676], bl[9677], bl[9678], bl[9679], bl[9680], bl[9681], bl[9682], bl[9683], bl[9684], bl[9685], bl[9686], bl[9687], bl[9688], bl[9689], bl[9690], bl[9691], bl[9692], bl[9693], bl[9694], bl[9695], bl[9696], bl[9697], bl[9698], bl[9699], bl[9700], bl[9701], bl[9702], bl[9703], bl[9704], bl[9705], bl[9706], bl[9707], bl[9708], bl[9709], bl[9710], bl[9711], bl[9712], bl[9713], bl[9714], bl[9715], bl[9716], bl[9717], bl[9718], bl[9719], bl[9720], bl[9721], bl[9722], bl[9723], bl[9724], bl[9725], bl[9726], bl[9727], bl[9728], bl[9729], bl[9730], bl[9731], bl[9732], bl[9733], bl[9734], bl[9735], bl[9736], bl[9737], bl[9738], bl[9739], bl[9740], bl[9741], bl[9742], bl[9743], bl[9744], bl[9745], bl[9746], bl[9747], bl[9748], bl[9749], bl[9750], bl[9751], bl[9752], bl[9753], bl[9754], bl[9755], bl[9756], bl[9757], bl[9758], bl[9759], bl[9760], bl[9761], bl[9762], bl[9763], bl[9764], bl[9765], bl[9766], bl[9767], bl[9768], bl[9769], bl[9770], bl[9771], bl[9772], bl[9773], bl[9774], bl[9775], bl[9776], bl[9777], bl[9778], bl[9779], bl[9780], bl[9781], bl[9782], bl[9783], bl[9784], bl[9785], bl[9786], bl[9787], bl[9788], bl[9789], bl[9790], bl[9791], bl[9792], bl[9793], bl[9794], bl[9795], bl[9796], bl[9797], bl[9798], bl[9799], bl[9800], bl[9801], bl[9802], bl[9803], bl[9804], bl[9805], bl[9806], bl[9807], bl[9808], bl[9809], bl[9810], bl[9811], bl[9812], bl[9813], bl[9814], bl[9815], bl[9816], bl[9817], bl[9818], bl[9819], bl[9820], bl[9821], bl[9822], bl[9823], bl[9824], bl[9825], bl[9826], bl[9827], bl[9828], bl[9829], bl[9830], bl[9831], bl[9832], bl[9833], bl[9834], bl[9835], bl[9836], bl[9837], bl[9838], bl[9839], bl[9840], bl[9841], bl[9842], bl[9843], bl[9844], bl[9845], bl[9846], bl[9847], bl[9848], bl[9849], bl[9850], bl[9851], bl[9852], bl[9853], bl[9854], bl[9855], bl[9856], bl[9857], bl[9858], bl[9859], bl[9860], bl[9861], bl[9862], bl[9863], bl[9864], bl[9865], bl[9866], bl[9867], bl[9868], bl[9869], bl[9870], bl[9871], bl[9872], bl[9873], bl[9874], bl[9875], bl[9876], bl[9877], bl[9878], bl[9879], bl[9880], bl[9881], bl[9882], bl[9883], bl[9884], bl[9885], bl[9886], bl[9887], bl[9888], bl[9889], bl[9890], bl[9891], bl[9892], bl[9893], bl[9894], bl[9895], bl[9896], bl[9897], bl[9898], bl[9899], bl[9900], bl[9901], bl[9902], bl[9903], bl[9904], bl[9905], bl[9906], bl[9907], bl[9908], bl[9909], bl[9910], bl[9911], bl[9912], bl[9913], bl[9914], bl[9915], bl[9916], bl[9917], bl[9918], bl[9919], bl[9920], bl[9921], bl[9922], bl[9923], bl[9924], bl[9925], bl[9926], bl[9927], bl[9928], bl[9929], bl[9930], bl[9931], bl[9932], bl[9933], bl[9934], bl[9935], bl[9936], bl[9937], bl[9938], bl[9939], bl[9940], bl[9941], bl[9942], bl[9943], bl[9944], bl[9945], bl[9946], bl[9947], bl[9948], bl[9949], bl[9950], bl[9951], bl[9952], bl[9953], bl[9954], bl[9955], bl[9956], bl[9957], bl[9958], bl[9959], bl[9960], bl[9961], bl[9962], bl[9963], bl[9964], bl[9965], bl[9966], bl[9967], bl[9968], bl[9969], bl[9970], bl[9971], bl[9972], bl[9973], bl[9974], bl[9975], bl[9976], bl[9977], bl[9978], bl[9979], bl[9980], bl[9981], bl[9982], bl[9983], bl[9984], bl[9985], bl[9986], bl[9987], bl[9988], bl[9989], bl[9990], bl[9991], bl[9992], bl[9993], bl[9994], bl[9995], bl[9996], bl[9997], bl[9998], bl[9999], bl[10000], bl[10001], bl[10002], bl[10003], bl[10004], bl[10005], bl[10006], bl[10007], bl[10008], bl[10009], bl[10010], bl[10011], bl[10012], bl[10013], bl[10014], bl[10015], bl[10016], bl[10017], bl[10018], bl[10019], bl[10020], bl[10021], bl[10022], bl[10023], bl[10024], bl[10025], bl[10026], bl[10027], bl[10028], bl[10029], bl[10030], bl[10031], bl[10032], bl[10033], bl[10034], bl[10035], bl[10036], bl[10037], bl[10038], bl[10039], bl[10040], bl[10041], bl[10042], bl[10043], bl[10044], bl[10045], bl[10046], bl[10047], bl[10048], bl[10049], bl[10050], bl[10051], bl[10052], bl[10053], bl[10054], bl[10055], bl[10056], bl[10057], bl[10058], bl[10059], bl[10060], bl[10061], bl[10062], bl[10063], bl[10064], bl[10065], bl[10066], bl[10067], bl[10068], bl[10069], bl[10070], bl[10071], bl[10072], bl[10073], bl[10074], bl[10075], bl[10076], bl[10077], bl[10078], bl[10079], bl[10080], bl[10081], bl[10082], bl[10083], bl[10084], bl[10085], bl[10086], bl[10087], bl[10088], bl[10089], bl[10090], bl[10091], bl[10092], bl[10093], bl[10094], bl[10095], bl[10096], bl[10097], bl[10098], bl[10099], bl[10100], bl[10101], bl[10102], bl[10103], bl[10104], bl[10105], bl[10106], bl[10107], bl[10108], bl[10109], bl[10110], bl[10111], bl[10112], bl[10113], bl[10114], bl[10115], bl[10116], bl[10117], bl[10118], bl[10119], bl[10120], bl[10121], bl[10122], bl[10123], bl[10124], bl[10125], bl[10126], bl[10127], bl[10128], bl[10129], bl[10130], bl[10131], bl[10132], bl[10133], bl[10134], bl[10135], bl[10136], bl[10137], bl[10138], bl[10139], bl[10140], bl[10141], bl[10142], bl[10143], bl[10144], bl[10145], bl[10146], bl[10147], bl[10148], bl[10149], bl[10150], bl[10151], bl[10152], bl[10153], bl[10154], bl[10155], bl[10156], bl[10157], bl[10158], bl[10159], bl[10160], bl[10161], bl[10162], bl[10163], bl[10164], bl[10165], bl[10166], bl[10167], bl[10168], bl[10169], bl[10170], bl[10171], bl[10172], bl[10173], bl[10174], bl[10175], bl[10176], bl[10177], bl[10178], bl[10179], bl[10180], bl[10181], bl[10182], bl[10183], bl[12784], bl[12785], bl[12786], bl[12787], bl[12788], bl[12789], bl[12790], bl[12791], bl[12792], bl[12793], bl[12794], bl[12795], bl[12796], bl[12797], bl[12798], bl[12799], bl[12800], bl[12801], bl[12802], bl[12803], bl[12804], bl[12805], bl[12806], bl[12807], bl[12808], bl[12809], bl[12810], bl[12811], bl[12812], bl[12813], bl[12814], bl[12815], bl[12816], bl[12817], bl[12818], bl[12819], bl[12820], bl[12821], bl[12822], bl[12823], bl[12824], bl[12825], bl[12826], bl[12827], bl[12828], bl[12829], bl[12830], bl[12831], bl[12832], bl[12833], bl[12834], bl[12835], bl[12836], bl[12837], bl[12838], bl[12839], bl[12840], bl[12841], bl[12842], bl[12843], bl[12844], bl[12845], bl[12846], bl[12847], bl[12848], bl[12849], bl[12850], bl[12851], bl[12852], bl[12853], bl[12854], bl[12855], bl[12856], bl[12857], bl[12858], bl[12859], bl[12860], bl[12861], bl[12862], bl[12863], bl[9084], bl[9085], bl[9086], bl[9087], bl[9088], bl[9089], bl[9090], bl[9091], bl[9092], bl[9093], bl[9094], bl[9095], bl[9096], bl[9097], bl[9098], bl[9099], bl[9100], bl[9101], bl[9102], bl[9103], bl[9104], bl[9105], bl[9106], bl[9107], bl[9108], bl[9109], bl[9110], bl[9111], bl[9112], bl[9113], bl[9114], bl[9115], bl[9116], bl[9117], bl[9118], bl[9119], bl[9120], bl[9121], bl[9122], bl[9123], bl[9124], bl[9125], bl[9126], bl[9127], bl[9128], bl[9129], bl[9130], bl[9131], bl[9132], bl[9133], bl[9134], bl[9135], bl[9136], bl[9137], bl[9138], bl[9139], bl[9140], bl[9141], bl[9142], bl[9143], bl[9144], bl[9145], bl[9146], bl[9147], bl[9148], bl[9149], bl[9150], bl[9151], bl[9152], bl[9153], bl[9154], bl[9155], bl[9156], bl[9157], bl[9158], bl[9159], bl[9160], bl[9161], bl[9162], bl[9163], bl[12704], bl[12705], bl[12706], bl[12707], bl[12708], bl[12709], bl[12710], bl[12711], bl[12712], bl[12713], bl[12714], bl[12715], bl[12716], bl[12717], bl[12718], bl[12719], bl[12720], bl[12721], bl[12722], bl[12723], bl[12724], bl[12725], bl[12726], bl[12727], bl[12728], bl[12729], bl[12730], bl[12731], bl[12732], bl[12733], bl[12734], bl[12735], bl[12736], bl[12737], bl[12738], bl[12739], bl[12740], bl[12741], bl[12742], bl[12743], bl[12744], bl[12745], bl[12746], bl[12747], bl[12748], bl[12749], bl[12750], bl[12751], bl[12752], bl[12753], bl[12754], bl[12755], bl[12756], bl[12757], bl[12758], bl[12759], bl[12760], bl[12761], bl[12762], bl[12763], bl[12764], bl[12765], bl[12766], bl[12767], bl[12768], bl[12769], bl[12770], bl[12771], bl[12772], bl[12773], bl[12774], bl[12775], bl[12776], bl[12777], bl[12778], bl[12779], bl[12780], bl[12781], bl[12782], bl[12783]}),
        .wl({wl[9164], wl[9165], wl[9166], wl[9167], wl[9168], wl[9169], wl[9170], wl[9171], wl[9172], wl[9173], wl[9174], wl[9175], wl[9176], wl[9177], wl[9178], wl[9179], wl[9180], wl[9181], wl[9182], wl[9183], wl[9184], wl[9185], wl[9186], wl[9187], wl[9188], wl[9189], wl[9190], wl[9191], wl[9192], wl[9193], wl[9194], wl[9195], wl[9196], wl[9197], wl[9198], wl[9199], wl[9200], wl[9201], wl[9202], wl[9203], wl[9204], wl[9205], wl[9206], wl[9207], wl[9208], wl[9209], wl[9210], wl[9211], wl[9212], wl[9213], wl[9214], wl[9215], wl[9216], wl[9217], wl[9218], wl[9219], wl[9220], wl[9221], wl[9222], wl[9223], wl[9224], wl[9225], wl[9226], wl[9227], wl[9228], wl[9229], wl[9230], wl[9231], wl[9232], wl[9233], wl[9234], wl[9235], wl[9236], wl[9237], wl[9238], wl[9239], wl[9240], wl[9241], wl[9242], wl[9243], wl[9244], wl[9245], wl[9246], wl[9247], wl[9248], wl[9249], wl[9250], wl[9251], wl[9252], wl[9253], wl[9254], wl[9255], wl[9256], wl[9257], wl[9258], wl[9259], wl[9260], wl[9261], wl[9262], wl[9263], wl[9264], wl[9265], wl[9266], wl[9267], wl[9268], wl[9269], wl[9270], wl[9271], wl[9272], wl[9273], wl[9274], wl[9275], wl[9276], wl[9277], wl[9278], wl[9279], wl[9280], wl[9281], wl[9282], wl[9283], wl[9284], wl[9285], wl[9286], wl[9287], wl[9288], wl[9289], wl[9290], wl[9291], wl[9292], wl[9293], wl[9294], wl[9295], wl[9296], wl[9297], wl[9298], wl[9299], wl[9300], wl[9301], wl[9302], wl[9303], wl[9304], wl[9305], wl[9306], wl[9307], wl[9308], wl[9309], wl[9310], wl[9311], wl[9312], wl[9313], wl[9314], wl[9315], wl[9316], wl[9317], wl[9318], wl[9319], wl[9320], wl[9321], wl[9322], wl[9323], wl[9324], wl[9325], wl[9326], wl[9327], wl[9328], wl[9329], wl[9330], wl[9331], wl[9332], wl[9333], wl[9334], wl[9335], wl[9336], wl[9337], wl[9338], wl[9339], wl[9340], wl[9341], wl[9342], wl[9343], wl[9344], wl[9345], wl[9346], wl[9347], wl[9348], wl[9349], wl[9350], wl[9351], wl[9352], wl[9353], wl[9354], wl[9355], wl[9356], wl[9357], wl[9358], wl[9359], wl[9360], wl[9361], wl[9362], wl[9363], wl[9364], wl[9365], wl[9366], wl[9367], wl[9368], wl[9369], wl[9370], wl[9371], wl[9372], wl[9373], wl[9374], wl[9375], wl[9376], wl[9377], wl[9378], wl[9379], wl[9380], wl[9381], wl[9382], wl[9383], wl[9384], wl[9385], wl[9386], wl[9387], wl[9388], wl[9389], wl[9390], wl[9391], wl[9392], wl[9393], wl[9394], wl[9395], wl[9396], wl[9397], wl[9398], wl[9399], wl[9400], wl[9401], wl[9402], wl[9403], wl[9404], wl[9405], wl[9406], wl[9407], wl[9408], wl[9409], wl[9410], wl[9411], wl[9412], wl[9413], wl[9414], wl[9415], wl[9416], wl[9417], wl[9418], wl[9419], wl[9420], wl[9421], wl[9422], wl[9423], wl[9424], wl[9425], wl[9426], wl[9427], wl[9428], wl[9429], wl[9430], wl[9431], wl[9432], wl[9433], wl[9434], wl[9435], wl[9436], wl[9437], wl[9438], wl[9439], wl[9440], wl[9441], wl[9442], wl[9443], wl[9444], wl[9445], wl[9446], wl[9447], wl[9448], wl[9449], wl[9450], wl[9451], wl[9452], wl[9453], wl[9454], wl[9455], wl[9456], wl[9457], wl[9458], wl[9459], wl[9460], wl[9461], wl[9462], wl[9463], wl[9464], wl[9465], wl[9466], wl[9467], wl[9468], wl[9469], wl[9470], wl[9471], wl[9472], wl[9473], wl[9474], wl[9475], wl[9476], wl[9477], wl[9478], wl[9479], wl[9480], wl[9481], wl[9482], wl[9483], wl[9484], wl[9485], wl[9486], wl[9487], wl[9488], wl[9489], wl[9490], wl[9491], wl[9492], wl[9493], wl[9494], wl[9495], wl[9496], wl[9497], wl[9498], wl[9499], wl[9500], wl[9501], wl[9502], wl[9503], wl[9504], wl[9505], wl[9506], wl[9507], wl[9508], wl[9509], wl[9510], wl[9511], wl[9512], wl[9513], wl[9514], wl[9515], wl[9516], wl[9517], wl[9518], wl[9519], wl[9520], wl[9521], wl[9522], wl[9523], wl[9524], wl[9525], wl[9526], wl[9527], wl[9528], wl[9529], wl[9530], wl[9531], wl[9532], wl[9533], wl[9534], wl[9535], wl[9536], wl[9537], wl[9538], wl[9539], wl[9540], wl[9541], wl[9542], wl[9543], wl[9544], wl[9545], wl[9546], wl[9547], wl[9548], wl[9549], wl[9550], wl[9551], wl[9552], wl[9553], wl[9554], wl[9555], wl[9556], wl[9557], wl[9558], wl[9559], wl[9560], wl[9561], wl[9562], wl[9563], wl[9564], wl[9565], wl[9566], wl[9567], wl[9568], wl[9569], wl[9570], wl[9571], wl[9572], wl[9573], wl[9574], wl[9575], wl[9576], wl[9577], wl[9578], wl[9579], wl[9580], wl[9581], wl[9582], wl[9583], wl[9584], wl[9585], wl[9586], wl[9587], wl[9588], wl[9589], wl[9590], wl[9591], wl[9592], wl[9593], wl[9594], wl[9595], wl[9596], wl[9597], wl[9598], wl[9599], wl[9600], wl[9601], wl[9602], wl[9603], wl[9604], wl[9605], wl[9606], wl[9607], wl[9608], wl[9609], wl[9610], wl[9611], wl[9612], wl[9613], wl[9614], wl[9615], wl[9616], wl[9617], wl[9618], wl[9619], wl[9620], wl[9621], wl[9622], wl[9623], wl[9624], wl[9625], wl[9626], wl[9627], wl[9628], wl[9629], wl[9630], wl[9631], wl[9632], wl[9633], wl[9634], wl[9635], wl[9636], wl[9637], wl[9638], wl[9639], wl[9640], wl[9641], wl[9642], wl[9643], wl[9644], wl[9645], wl[9646], wl[9647], wl[9648], wl[9649], wl[9650], wl[9651], wl[9652], wl[9653], wl[9654], wl[9655], wl[9656], wl[9657], wl[9658], wl[9659], wl[9660], wl[9661], wl[9662], wl[9663], wl[9664], wl[9665], wl[9666], wl[9667], wl[9668], wl[9669], wl[9670], wl[9671], wl[9672], wl[9673], wl[9674], wl[9675], wl[9676], wl[9677], wl[9678], wl[9679], wl[9680], wl[9681], wl[9682], wl[9683], wl[9684], wl[9685], wl[9686], wl[9687], wl[9688], wl[9689], wl[9690], wl[9691], wl[9692], wl[9693], wl[9694], wl[9695], wl[9696], wl[9697], wl[9698], wl[9699], wl[9700], wl[9701], wl[9702], wl[9703], wl[9704], wl[9705], wl[9706], wl[9707], wl[9708], wl[9709], wl[9710], wl[9711], wl[9712], wl[9713], wl[9714], wl[9715], wl[9716], wl[9717], wl[9718], wl[9719], wl[9720], wl[9721], wl[9722], wl[9723], wl[9724], wl[9725], wl[9726], wl[9727], wl[9728], wl[9729], wl[9730], wl[9731], wl[9732], wl[9733], wl[9734], wl[9735], wl[9736], wl[9737], wl[9738], wl[9739], wl[9740], wl[9741], wl[9742], wl[9743], wl[9744], wl[9745], wl[9746], wl[9747], wl[9748], wl[9749], wl[9750], wl[9751], wl[9752], wl[9753], wl[9754], wl[9755], wl[9756], wl[9757], wl[9758], wl[9759], wl[9760], wl[9761], wl[9762], wl[9763], wl[9764], wl[9765], wl[9766], wl[9767], wl[9768], wl[9769], wl[9770], wl[9771], wl[9772], wl[9773], wl[9774], wl[9775], wl[9776], wl[9777], wl[9778], wl[9779], wl[9780], wl[9781], wl[9782], wl[9783], wl[9784], wl[9785], wl[9786], wl[9787], wl[9788], wl[9789], wl[9790], wl[9791], wl[9792], wl[9793], wl[9794], wl[9795], wl[9796], wl[9797], wl[9798], wl[9799], wl[9800], wl[9801], wl[9802], wl[9803], wl[9804], wl[9805], wl[9806], wl[9807], wl[9808], wl[9809], wl[9810], wl[9811], wl[9812], wl[9813], wl[9814], wl[9815], wl[9816], wl[9817], wl[9818], wl[9819], wl[9820], wl[9821], wl[9822], wl[9823], wl[9824], wl[9825], wl[9826], wl[9827], wl[9828], wl[9829], wl[9830], wl[9831], wl[9832], wl[9833], wl[9834], wl[9835], wl[9836], wl[9837], wl[9838], wl[9839], wl[9840], wl[9841], wl[9842], wl[9843], wl[9844], wl[9845], wl[9846], wl[9847], wl[9848], wl[9849], wl[9850], wl[9851], wl[9852], wl[9853], wl[9854], wl[9855], wl[9856], wl[9857], wl[9858], wl[9859], wl[9860], wl[9861], wl[9862], wl[9863], wl[9864], wl[9865], wl[9866], wl[9867], wl[9868], wl[9869], wl[9870], wl[9871], wl[9872], wl[9873], wl[9874], wl[9875], wl[9876], wl[9877], wl[9878], wl[9879], wl[9880], wl[9881], wl[9882], wl[9883], wl[9884], wl[9885], wl[9886], wl[9887], wl[9888], wl[9889], wl[9890], wl[9891], wl[9892], wl[9893], wl[9894], wl[9895], wl[9896], wl[9897], wl[9898], wl[9899], wl[9900], wl[9901], wl[9902], wl[9903], wl[9904], wl[9905], wl[9906], wl[9907], wl[9908], wl[9909], wl[9910], wl[9911], wl[9912], wl[9913], wl[9914], wl[9915], wl[9916], wl[9917], wl[9918], wl[9919], wl[9920], wl[9921], wl[9922], wl[9923], wl[9924], wl[9925], wl[9926], wl[9927], wl[9928], wl[9929], wl[9930], wl[9931], wl[9932], wl[9933], wl[9934], wl[9935], wl[9936], wl[9937], wl[9938], wl[9939], wl[9940], wl[9941], wl[9942], wl[9943], wl[9944], wl[9945], wl[9946], wl[9947], wl[9948], wl[9949], wl[9950], wl[9951], wl[9952], wl[9953], wl[9954], wl[9955], wl[9956], wl[9957], wl[9958], wl[9959], wl[9960], wl[9961], wl[9962], wl[9963], wl[9964], wl[9965], wl[9966], wl[9967], wl[9968], wl[9969], wl[9970], wl[9971], wl[9972], wl[9973], wl[9974], wl[9975], wl[9976], wl[9977], wl[9978], wl[9979], wl[9980], wl[9981], wl[9982], wl[9983], wl[9984], wl[9985], wl[9986], wl[9987], wl[9988], wl[9989], wl[9990], wl[9991], wl[9992], wl[9993], wl[9994], wl[9995], wl[9996], wl[9997], wl[9998], wl[9999], wl[10000], wl[10001], wl[10002], wl[10003], wl[10004], wl[10005], wl[10006], wl[10007], wl[10008], wl[10009], wl[10010], wl[10011], wl[10012], wl[10013], wl[10014], wl[10015], wl[10016], wl[10017], wl[10018], wl[10019], wl[10020], wl[10021], wl[10022], wl[10023], wl[10024], wl[10025], wl[10026], wl[10027], wl[10028], wl[10029], wl[10030], wl[10031], wl[10032], wl[10033], wl[10034], wl[10035], wl[10036], wl[10037], wl[10038], wl[10039], wl[10040], wl[10041], wl[10042], wl[10043], wl[10044], wl[10045], wl[10046], wl[10047], wl[10048], wl[10049], wl[10050], wl[10051], wl[10052], wl[10053], wl[10054], wl[10055], wl[10056], wl[10057], wl[10058], wl[10059], wl[10060], wl[10061], wl[10062], wl[10063], wl[10064], wl[10065], wl[10066], wl[10067], wl[10068], wl[10069], wl[10070], wl[10071], wl[10072], wl[10073], wl[10074], wl[10075], wl[10076], wl[10077], wl[10078], wl[10079], wl[10080], wl[10081], wl[10082], wl[10083], wl[10084], wl[10085], wl[10086], wl[10087], wl[10088], wl[10089], wl[10090], wl[10091], wl[10092], wl[10093], wl[10094], wl[10095], wl[10096], wl[10097], wl[10098], wl[10099], wl[10100], wl[10101], wl[10102], wl[10103], wl[10104], wl[10105], wl[10106], wl[10107], wl[10108], wl[10109], wl[10110], wl[10111], wl[10112], wl[10113], wl[10114], wl[10115], wl[10116], wl[10117], wl[10118], wl[10119], wl[10120], wl[10121], wl[10122], wl[10123], wl[10124], wl[10125], wl[10126], wl[10127], wl[10128], wl[10129], wl[10130], wl[10131], wl[10132], wl[10133], wl[10134], wl[10135], wl[10136], wl[10137], wl[10138], wl[10139], wl[10140], wl[10141], wl[10142], wl[10143], wl[10144], wl[10145], wl[10146], wl[10147], wl[10148], wl[10149], wl[10150], wl[10151], wl[10152], wl[10153], wl[10154], wl[10155], wl[10156], wl[10157], wl[10158], wl[10159], wl[10160], wl[10161], wl[10162], wl[10163], wl[10164], wl[10165], wl[10166], wl[10167], wl[10168], wl[10169], wl[10170], wl[10171], wl[10172], wl[10173], wl[10174], wl[10175], wl[10176], wl[10177], wl[10178], wl[10179], wl[10180], wl[10181], wl[10182], wl[10183], wl[12784], wl[12785], wl[12786], wl[12787], wl[12788], wl[12789], wl[12790], wl[12791], wl[12792], wl[12793], wl[12794], wl[12795], wl[12796], wl[12797], wl[12798], wl[12799], wl[12800], wl[12801], wl[12802], wl[12803], wl[12804], wl[12805], wl[12806], wl[12807], wl[12808], wl[12809], wl[12810], wl[12811], wl[12812], wl[12813], wl[12814], wl[12815], wl[12816], wl[12817], wl[12818], wl[12819], wl[12820], wl[12821], wl[12822], wl[12823], wl[12824], wl[12825], wl[12826], wl[12827], wl[12828], wl[12829], wl[12830], wl[12831], wl[12832], wl[12833], wl[12834], wl[12835], wl[12836], wl[12837], wl[12838], wl[12839], wl[12840], wl[12841], wl[12842], wl[12843], wl[12844], wl[12845], wl[12846], wl[12847], wl[12848], wl[12849], wl[12850], wl[12851], wl[12852], wl[12853], wl[12854], wl[12855], wl[12856], wl[12857], wl[12858], wl[12859], wl[12860], wl[12861], wl[12862], wl[12863], wl[9084], wl[9085], wl[9086], wl[9087], wl[9088], wl[9089], wl[9090], wl[9091], wl[9092], wl[9093], wl[9094], wl[9095], wl[9096], wl[9097], wl[9098], wl[9099], wl[9100], wl[9101], wl[9102], wl[9103], wl[9104], wl[9105], wl[9106], wl[9107], wl[9108], wl[9109], wl[9110], wl[9111], wl[9112], wl[9113], wl[9114], wl[9115], wl[9116], wl[9117], wl[9118], wl[9119], wl[9120], wl[9121], wl[9122], wl[9123], wl[9124], wl[9125], wl[9126], wl[9127], wl[9128], wl[9129], wl[9130], wl[9131], wl[9132], wl[9133], wl[9134], wl[9135], wl[9136], wl[9137], wl[9138], wl[9139], wl[9140], wl[9141], wl[9142], wl[9143], wl[9144], wl[9145], wl[9146], wl[9147], wl[9148], wl[9149], wl[9150], wl[9151], wl[9152], wl[9153], wl[9154], wl[9155], wl[9156], wl[9157], wl[9158], wl[9159], wl[9160], wl[9161], wl[9162], wl[9163], wl[12704], wl[12705], wl[12706], wl[12707], wl[12708], wl[12709], wl[12710], wl[12711], wl[12712], wl[12713], wl[12714], wl[12715], wl[12716], wl[12717], wl[12718], wl[12719], wl[12720], wl[12721], wl[12722], wl[12723], wl[12724], wl[12725], wl[12726], wl[12727], wl[12728], wl[12729], wl[12730], wl[12731], wl[12732], wl[12733], wl[12734], wl[12735], wl[12736], wl[12737], wl[12738], wl[12739], wl[12740], wl[12741], wl[12742], wl[12743], wl[12744], wl[12745], wl[12746], wl[12747], wl[12748], wl[12749], wl[12750], wl[12751], wl[12752], wl[12753], wl[12754], wl[12755], wl[12756], wl[12757], wl[12758], wl[12759], wl[12760], wl[12761], wl[12762], wl[12763], wl[12764], wl[12765], wl[12766], wl[12767], wl[12768], wl[12769], wl[12770], wl[12771], wl[12772], wl[12773], wl[12774], wl[12775], wl[12776], wl[12777], wl[12778], wl[12779], wl[12780], wl[12781], wl[12782], wl[12783]})
    );
    tile tile_3__4_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_1__3__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_1__3__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_1__3__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_2__2__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_2__2__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_2__2__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_1__2__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_1__2__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_1__2__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_1__2__grid_top_r_in[1]),
        .grid_left_in(grid_clb_2__3__grid_left_in),
        .grid_bottom_in(grid_clb_2__3__grid_bottom_in),
        .chanx_left_in(sb_1__1__2_chanx_right_out),
        .chanx_left_out(cbx_1__1__5_chanx_left_out),
        .grid_top_out(grid_clb_2__4__grid_bottom_in),
        .chany_bottom_in(sb_1__1__4_chany_top_out),
        .chany_bottom_out(cby_1__1__6_chany_bottom_out),
        .grid_right_out(grid_clb_3__3__grid_left_in),
        .chany_top_in_0(cby_1__1__7_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__8_chanx_left_out),
        .chany_top_out_0(sb_1__1__5_chany_top_out),
        .chanx_right_out_0(sb_1__1__5_chanx_right_out),
        .grid_top_r_in(sb_2__3__grid_top_r_in),
        .grid_top_l_in(sb_2__3__grid_top_l_in),
        .grid_right_t_in(sb_2__3__grid_right_t_in),
        .grid_right_b_in(sb_2__3__grid_right_b_in),
        .grid_bottom_r_in(sb_2__2__grid_top_r_in),
        .grid_bottom_l_in(sb_2__2__grid_top_l_in),
        .grid_left_t_in(sb_1__3__grid_right_t_in),
        .grid_left_b_in(sb_1__3__grid_right_b_in),
        .bl({bl[12944], bl[12945], bl[12946], bl[12947], bl[12948], bl[12949], bl[12950], bl[12951], bl[12952], bl[12953], bl[12954], bl[12955], bl[12956], bl[12957], bl[12958], bl[12959], bl[12960], bl[12961], bl[12962], bl[12963], bl[12964], bl[12965], bl[12966], bl[12967], bl[12968], bl[12969], bl[12970], bl[12971], bl[12972], bl[12973], bl[12974], bl[12975], bl[12976], bl[12977], bl[12978], bl[12979], bl[12980], bl[12981], bl[12982], bl[12983], bl[12984], bl[12985], bl[12986], bl[12987], bl[12988], bl[12989], bl[12990], bl[12991], bl[12992], bl[12993], bl[12994], bl[12995], bl[12996], bl[12997], bl[12998], bl[12999], bl[13000], bl[13001], bl[13002], bl[13003], bl[13004], bl[13005], bl[13006], bl[13007], bl[13008], bl[13009], bl[13010], bl[13011], bl[13012], bl[13013], bl[13014], bl[13015], bl[13016], bl[13017], bl[13018], bl[13019], bl[13020], bl[13021], bl[13022], bl[13023], bl[13024], bl[13025], bl[13026], bl[13027], bl[13028], bl[13029], bl[13030], bl[13031], bl[13032], bl[13033], bl[13034], bl[13035], bl[13036], bl[13037], bl[13038], bl[13039], bl[13040], bl[13041], bl[13042], bl[13043], bl[13044], bl[13045], bl[13046], bl[13047], bl[13048], bl[13049], bl[13050], bl[13051], bl[13052], bl[13053], bl[13054], bl[13055], bl[13056], bl[13057], bl[13058], bl[13059], bl[13060], bl[13061], bl[13062], bl[13063], bl[13064], bl[13065], bl[13066], bl[13067], bl[13068], bl[13069], bl[13070], bl[13071], bl[13072], bl[13073], bl[13074], bl[13075], bl[13076], bl[13077], bl[13078], bl[13079], bl[13080], bl[13081], bl[13082], bl[13083], bl[13084], bl[13085], bl[13086], bl[13087], bl[13088], bl[13089], bl[13090], bl[13091], bl[13092], bl[13093], bl[13094], bl[13095], bl[13096], bl[13097], bl[13098], bl[13099], bl[13100], bl[13101], bl[13102], bl[13103], bl[13104], bl[13105], bl[13106], bl[13107], bl[13108], bl[13109], bl[13110], bl[13111], bl[13112], bl[13113], bl[13114], bl[13115], bl[13116], bl[13117], bl[13118], bl[13119], bl[13120], bl[13121], bl[13122], bl[13123], bl[13124], bl[13125], bl[13126], bl[13127], bl[13128], bl[13129], bl[13130], bl[13131], bl[13132], bl[13133], bl[13134], bl[13135], bl[13136], bl[13137], bl[13138], bl[13139], bl[13140], bl[13141], bl[13142], bl[13143], bl[13144], bl[13145], bl[13146], bl[13147], bl[13148], bl[13149], bl[13150], bl[13151], bl[13152], bl[13153], bl[13154], bl[13155], bl[13156], bl[13157], bl[13158], bl[13159], bl[13160], bl[13161], bl[13162], bl[13163], bl[13164], bl[13165], bl[13166], bl[13167], bl[13168], bl[13169], bl[13170], bl[13171], bl[13172], bl[13173], bl[13174], bl[13175], bl[13176], bl[13177], bl[13178], bl[13179], bl[13180], bl[13181], bl[13182], bl[13183], bl[13184], bl[13185], bl[13186], bl[13187], bl[13188], bl[13189], bl[13190], bl[13191], bl[13192], bl[13193], bl[13194], bl[13195], bl[13196], bl[13197], bl[13198], bl[13199], bl[13200], bl[13201], bl[13202], bl[13203], bl[13204], bl[13205], bl[13206], bl[13207], bl[13208], bl[13209], bl[13210], bl[13211], bl[13212], bl[13213], bl[13214], bl[13215], bl[13216], bl[13217], bl[13218], bl[13219], bl[13220], bl[13221], bl[13222], bl[13223], bl[13224], bl[13225], bl[13226], bl[13227], bl[13228], bl[13229], bl[13230], bl[13231], bl[13232], bl[13233], bl[13234], bl[13235], bl[13236], bl[13237], bl[13238], bl[13239], bl[13240], bl[13241], bl[13242], bl[13243], bl[13244], bl[13245], bl[13246], bl[13247], bl[13248], bl[13249], bl[13250], bl[13251], bl[13252], bl[13253], bl[13254], bl[13255], bl[13256], bl[13257], bl[13258], bl[13259], bl[13260], bl[13261], bl[13262], bl[13263], bl[13264], bl[13265], bl[13266], bl[13267], bl[13268], bl[13269], bl[13270], bl[13271], bl[13272], bl[13273], bl[13274], bl[13275], bl[13276], bl[13277], bl[13278], bl[13279], bl[13280], bl[13281], bl[13282], bl[13283], bl[13284], bl[13285], bl[13286], bl[13287], bl[13288], bl[13289], bl[13290], bl[13291], bl[13292], bl[13293], bl[13294], bl[13295], bl[13296], bl[13297], bl[13298], bl[13299], bl[13300], bl[13301], bl[13302], bl[13303], bl[13304], bl[13305], bl[13306], bl[13307], bl[13308], bl[13309], bl[13310], bl[13311], bl[13312], bl[13313], bl[13314], bl[13315], bl[13316], bl[13317], bl[13318], bl[13319], bl[13320], bl[13321], bl[13322], bl[13323], bl[13324], bl[13325], bl[13326], bl[13327], bl[13328], bl[13329], bl[13330], bl[13331], bl[13332], bl[13333], bl[13334], bl[13335], bl[13336], bl[13337], bl[13338], bl[13339], bl[13340], bl[13341], bl[13342], bl[13343], bl[13344], bl[13345], bl[13346], bl[13347], bl[13348], bl[13349], bl[13350], bl[13351], bl[13352], bl[13353], bl[13354], bl[13355], bl[13356], bl[13357], bl[13358], bl[13359], bl[13360], bl[13361], bl[13362], bl[13363], bl[13364], bl[13365], bl[13366], bl[13367], bl[13368], bl[13369], bl[13370], bl[13371], bl[13372], bl[13373], bl[13374], bl[13375], bl[13376], bl[13377], bl[13378], bl[13379], bl[13380], bl[13381], bl[13382], bl[13383], bl[13384], bl[13385], bl[13386], bl[13387], bl[13388], bl[13389], bl[13390], bl[13391], bl[13392], bl[13393], bl[13394], bl[13395], bl[13396], bl[13397], bl[13398], bl[13399], bl[13400], bl[13401], bl[13402], bl[13403], bl[13404], bl[13405], bl[13406], bl[13407], bl[13408], bl[13409], bl[13410], bl[13411], bl[13412], bl[13413], bl[13414], bl[13415], bl[13416], bl[13417], bl[13418], bl[13419], bl[13420], bl[13421], bl[13422], bl[13423], bl[13424], bl[13425], bl[13426], bl[13427], bl[13428], bl[13429], bl[13430], bl[13431], bl[13432], bl[13433], bl[13434], bl[13435], bl[13436], bl[13437], bl[13438], bl[13439], bl[13440], bl[13441], bl[13442], bl[13443], bl[13444], bl[13445], bl[13446], bl[13447], bl[13448], bl[13449], bl[13450], bl[13451], bl[13452], bl[13453], bl[13454], bl[13455], bl[13456], bl[13457], bl[13458], bl[13459], bl[13460], bl[13461], bl[13462], bl[13463], bl[13464], bl[13465], bl[13466], bl[13467], bl[13468], bl[13469], bl[13470], bl[13471], bl[13472], bl[13473], bl[13474], bl[13475], bl[13476], bl[13477], bl[13478], bl[13479], bl[13480], bl[13481], bl[13482], bl[13483], bl[13484], bl[13485], bl[13486], bl[13487], bl[13488], bl[13489], bl[13490], bl[13491], bl[13492], bl[13493], bl[13494], bl[13495], bl[13496], bl[13497], bl[13498], bl[13499], bl[13500], bl[13501], bl[13502], bl[13503], bl[13504], bl[13505], bl[13506], bl[13507], bl[13508], bl[13509], bl[13510], bl[13511], bl[13512], bl[13513], bl[13514], bl[13515], bl[13516], bl[13517], bl[13518], bl[13519], bl[13520], bl[13521], bl[13522], bl[13523], bl[13524], bl[13525], bl[13526], bl[13527], bl[13528], bl[13529], bl[13530], bl[13531], bl[13532], bl[13533], bl[13534], bl[13535], bl[13536], bl[13537], bl[13538], bl[13539], bl[13540], bl[13541], bl[13542], bl[13543], bl[13544], bl[13545], bl[13546], bl[13547], bl[13548], bl[13549], bl[13550], bl[13551], bl[13552], bl[13553], bl[13554], bl[13555], bl[13556], bl[13557], bl[13558], bl[13559], bl[13560], bl[13561], bl[13562], bl[13563], bl[13564], bl[13565], bl[13566], bl[13567], bl[13568], bl[13569], bl[13570], bl[13571], bl[13572], bl[13573], bl[13574], bl[13575], bl[13576], bl[13577], bl[13578], bl[13579], bl[13580], bl[13581], bl[13582], bl[13583], bl[13584], bl[13585], bl[13586], bl[13587], bl[13588], bl[13589], bl[13590], bl[13591], bl[13592], bl[13593], bl[13594], bl[13595], bl[13596], bl[13597], bl[13598], bl[13599], bl[13600], bl[13601], bl[13602], bl[13603], bl[13604], bl[13605], bl[13606], bl[13607], bl[13608], bl[13609], bl[13610], bl[13611], bl[13612], bl[13613], bl[13614], bl[13615], bl[13616], bl[13617], bl[13618], bl[13619], bl[13620], bl[13621], bl[13622], bl[13623], bl[13624], bl[13625], bl[13626], bl[13627], bl[13628], bl[13629], bl[13630], bl[13631], bl[13632], bl[13633], bl[13634], bl[13635], bl[13636], bl[13637], bl[13638], bl[13639], bl[13640], bl[13641], bl[13642], bl[13643], bl[13644], bl[13645], bl[13646], bl[13647], bl[13648], bl[13649], bl[13650], bl[13651], bl[13652], bl[13653], bl[13654], bl[13655], bl[13656], bl[13657], bl[13658], bl[13659], bl[13660], bl[13661], bl[13662], bl[13663], bl[13664], bl[13665], bl[13666], bl[13667], bl[13668], bl[13669], bl[13670], bl[13671], bl[13672], bl[13673], bl[13674], bl[13675], bl[13676], bl[13677], bl[13678], bl[13679], bl[13680], bl[13681], bl[13682], bl[13683], bl[13684], bl[13685], bl[13686], bl[13687], bl[13688], bl[13689], bl[13690], bl[13691], bl[13692], bl[13693], bl[13694], bl[13695], bl[13696], bl[13697], bl[13698], bl[13699], bl[13700], bl[13701], bl[13702], bl[13703], bl[13704], bl[13705], bl[13706], bl[13707], bl[13708], bl[13709], bl[13710], bl[13711], bl[13712], bl[13713], bl[13714], bl[13715], bl[13716], bl[13717], bl[13718], bl[13719], bl[13720], bl[13721], bl[13722], bl[13723], bl[13724], bl[13725], bl[13726], bl[13727], bl[13728], bl[13729], bl[13730], bl[13731], bl[13732], bl[13733], bl[13734], bl[13735], bl[13736], bl[13737], bl[13738], bl[13739], bl[13740], bl[13741], bl[13742], bl[13743], bl[13744], bl[13745], bl[13746], bl[13747], bl[13748], bl[13749], bl[13750], bl[13751], bl[13752], bl[13753], bl[13754], bl[13755], bl[13756], bl[13757], bl[13758], bl[13759], bl[13760], bl[13761], bl[13762], bl[13763], bl[13764], bl[13765], bl[13766], bl[13767], bl[13768], bl[13769], bl[13770], bl[13771], bl[13772], bl[13773], bl[13774], bl[13775], bl[13776], bl[13777], bl[13778], bl[13779], bl[13780], bl[13781], bl[13782], bl[13783], bl[13784], bl[13785], bl[13786], bl[13787], bl[13788], bl[13789], bl[13790], bl[13791], bl[13792], bl[13793], bl[13794], bl[13795], bl[13796], bl[13797], bl[13798], bl[13799], bl[13800], bl[13801], bl[13802], bl[13803], bl[13804], bl[13805], bl[13806], bl[13807], bl[13808], bl[13809], bl[13810], bl[13811], bl[13812], bl[13813], bl[13814], bl[13815], bl[13816], bl[13817], bl[13818], bl[13819], bl[13820], bl[13821], bl[13822], bl[13823], bl[13824], bl[13825], bl[13826], bl[13827], bl[13828], bl[13829], bl[13830], bl[13831], bl[13832], bl[13833], bl[13834], bl[13835], bl[13836], bl[13837], bl[13838], bl[13839], bl[13840], bl[13841], bl[13842], bl[13843], bl[13844], bl[13845], bl[13846], bl[13847], bl[13848], bl[13849], bl[13850], bl[13851], bl[13852], bl[13853], bl[13854], bl[13855], bl[13856], bl[13857], bl[13858], bl[13859], bl[13860], bl[13861], bl[13862], bl[13863], bl[13864], bl[13865], bl[13866], bl[13867], bl[13868], bl[13869], bl[13870], bl[13871], bl[13872], bl[13873], bl[13874], bl[13875], bl[13876], bl[13877], bl[13878], bl[13879], bl[13880], bl[13881], bl[13882], bl[13883], bl[13884], bl[13885], bl[13886], bl[13887], bl[13888], bl[13889], bl[13890], bl[13891], bl[13892], bl[13893], bl[13894], bl[13895], bl[13896], bl[13897], bl[13898], bl[13899], bl[13900], bl[13901], bl[13902], bl[13903], bl[13904], bl[13905], bl[13906], bl[13907], bl[13908], bl[13909], bl[13910], bl[13911], bl[13912], bl[13913], bl[13914], bl[13915], bl[13916], bl[13917], bl[13918], bl[13919], bl[13920], bl[13921], bl[13922], bl[13923], bl[13924], bl[13925], bl[13926], bl[13927], bl[13928], bl[13929], bl[13930], bl[13931], bl[13932], bl[13933], bl[13934], bl[13935], bl[13936], bl[13937], bl[13938], bl[13939], bl[13940], bl[13941], bl[13942], bl[13943], bl[13944], bl[13945], bl[13946], bl[13947], bl[13948], bl[13949], bl[13950], bl[13951], bl[13952], bl[13953], bl[13954], bl[13955], bl[13956], bl[13957], bl[13958], bl[13959], bl[13960], bl[13961], bl[13962], bl[13963], bl[19068], bl[19069], bl[19070], bl[19071], bl[19072], bl[19073], bl[19074], bl[19075], bl[19076], bl[19077], bl[19078], bl[19079], bl[19080], bl[19081], bl[19082], bl[19083], bl[19084], bl[19085], bl[19086], bl[19087], bl[19088], bl[19089], bl[19090], bl[19091], bl[19092], bl[19093], bl[19094], bl[19095], bl[19096], bl[19097], bl[19098], bl[19099], bl[19100], bl[19101], bl[19102], bl[19103], bl[19104], bl[19105], bl[19106], bl[19107], bl[19108], bl[19109], bl[19110], bl[19111], bl[19112], bl[19113], bl[19114], bl[19115], bl[19116], bl[19117], bl[19118], bl[19119], bl[19120], bl[19121], bl[19122], bl[19123], bl[19124], bl[19125], bl[19126], bl[19127], bl[19128], bl[19129], bl[19130], bl[19131], bl[19132], bl[19133], bl[19134], bl[19135], bl[19136], bl[19137], bl[19138], bl[19139], bl[19140], bl[19141], bl[19142], bl[19143], bl[19144], bl[19145], bl[19146], bl[19147], bl[12864], bl[12865], bl[12866], bl[12867], bl[12868], bl[12869], bl[12870], bl[12871], bl[12872], bl[12873], bl[12874], bl[12875], bl[12876], bl[12877], bl[12878], bl[12879], bl[12880], bl[12881], bl[12882], bl[12883], bl[12884], bl[12885], bl[12886], bl[12887], bl[12888], bl[12889], bl[12890], bl[12891], bl[12892], bl[12893], bl[12894], bl[12895], bl[12896], bl[12897], bl[12898], bl[12899], bl[12900], bl[12901], bl[12902], bl[12903], bl[12904], bl[12905], bl[12906], bl[12907], bl[12908], bl[12909], bl[12910], bl[12911], bl[12912], bl[12913], bl[12914], bl[12915], bl[12916], bl[12917], bl[12918], bl[12919], bl[12920], bl[12921], bl[12922], bl[12923], bl[12924], bl[12925], bl[12926], bl[12927], bl[12928], bl[12929], bl[12930], bl[12931], bl[12932], bl[12933], bl[12934], bl[12935], bl[12936], bl[12937], bl[12938], bl[12939], bl[12940], bl[12941], bl[12942], bl[12943], bl[18988], bl[18989], bl[18990], bl[18991], bl[18992], bl[18993], bl[18994], bl[18995], bl[18996], bl[18997], bl[18998], bl[18999], bl[19000], bl[19001], bl[19002], bl[19003], bl[19004], bl[19005], bl[19006], bl[19007], bl[19008], bl[19009], bl[19010], bl[19011], bl[19012], bl[19013], bl[19014], bl[19015], bl[19016], bl[19017], bl[19018], bl[19019], bl[19020], bl[19021], bl[19022], bl[19023], bl[19024], bl[19025], bl[19026], bl[19027], bl[19028], bl[19029], bl[19030], bl[19031], bl[19032], bl[19033], bl[19034], bl[19035], bl[19036], bl[19037], bl[19038], bl[19039], bl[19040], bl[19041], bl[19042], bl[19043], bl[19044], bl[19045], bl[19046], bl[19047], bl[19048], bl[19049], bl[19050], bl[19051], bl[19052], bl[19053], bl[19054], bl[19055], bl[19056], bl[19057], bl[19058], bl[19059], bl[19060], bl[19061], bl[19062], bl[19063], bl[19064], bl[19065], bl[19066], bl[19067]}),
        .wl({wl[12944], wl[12945], wl[12946], wl[12947], wl[12948], wl[12949], wl[12950], wl[12951], wl[12952], wl[12953], wl[12954], wl[12955], wl[12956], wl[12957], wl[12958], wl[12959], wl[12960], wl[12961], wl[12962], wl[12963], wl[12964], wl[12965], wl[12966], wl[12967], wl[12968], wl[12969], wl[12970], wl[12971], wl[12972], wl[12973], wl[12974], wl[12975], wl[12976], wl[12977], wl[12978], wl[12979], wl[12980], wl[12981], wl[12982], wl[12983], wl[12984], wl[12985], wl[12986], wl[12987], wl[12988], wl[12989], wl[12990], wl[12991], wl[12992], wl[12993], wl[12994], wl[12995], wl[12996], wl[12997], wl[12998], wl[12999], wl[13000], wl[13001], wl[13002], wl[13003], wl[13004], wl[13005], wl[13006], wl[13007], wl[13008], wl[13009], wl[13010], wl[13011], wl[13012], wl[13013], wl[13014], wl[13015], wl[13016], wl[13017], wl[13018], wl[13019], wl[13020], wl[13021], wl[13022], wl[13023], wl[13024], wl[13025], wl[13026], wl[13027], wl[13028], wl[13029], wl[13030], wl[13031], wl[13032], wl[13033], wl[13034], wl[13035], wl[13036], wl[13037], wl[13038], wl[13039], wl[13040], wl[13041], wl[13042], wl[13043], wl[13044], wl[13045], wl[13046], wl[13047], wl[13048], wl[13049], wl[13050], wl[13051], wl[13052], wl[13053], wl[13054], wl[13055], wl[13056], wl[13057], wl[13058], wl[13059], wl[13060], wl[13061], wl[13062], wl[13063], wl[13064], wl[13065], wl[13066], wl[13067], wl[13068], wl[13069], wl[13070], wl[13071], wl[13072], wl[13073], wl[13074], wl[13075], wl[13076], wl[13077], wl[13078], wl[13079], wl[13080], wl[13081], wl[13082], wl[13083], wl[13084], wl[13085], wl[13086], wl[13087], wl[13088], wl[13089], wl[13090], wl[13091], wl[13092], wl[13093], wl[13094], wl[13095], wl[13096], wl[13097], wl[13098], wl[13099], wl[13100], wl[13101], wl[13102], wl[13103], wl[13104], wl[13105], wl[13106], wl[13107], wl[13108], wl[13109], wl[13110], wl[13111], wl[13112], wl[13113], wl[13114], wl[13115], wl[13116], wl[13117], wl[13118], wl[13119], wl[13120], wl[13121], wl[13122], wl[13123], wl[13124], wl[13125], wl[13126], wl[13127], wl[13128], wl[13129], wl[13130], wl[13131], wl[13132], wl[13133], wl[13134], wl[13135], wl[13136], wl[13137], wl[13138], wl[13139], wl[13140], wl[13141], wl[13142], wl[13143], wl[13144], wl[13145], wl[13146], wl[13147], wl[13148], wl[13149], wl[13150], wl[13151], wl[13152], wl[13153], wl[13154], wl[13155], wl[13156], wl[13157], wl[13158], wl[13159], wl[13160], wl[13161], wl[13162], wl[13163], wl[13164], wl[13165], wl[13166], wl[13167], wl[13168], wl[13169], wl[13170], wl[13171], wl[13172], wl[13173], wl[13174], wl[13175], wl[13176], wl[13177], wl[13178], wl[13179], wl[13180], wl[13181], wl[13182], wl[13183], wl[13184], wl[13185], wl[13186], wl[13187], wl[13188], wl[13189], wl[13190], wl[13191], wl[13192], wl[13193], wl[13194], wl[13195], wl[13196], wl[13197], wl[13198], wl[13199], wl[13200], wl[13201], wl[13202], wl[13203], wl[13204], wl[13205], wl[13206], wl[13207], wl[13208], wl[13209], wl[13210], wl[13211], wl[13212], wl[13213], wl[13214], wl[13215], wl[13216], wl[13217], wl[13218], wl[13219], wl[13220], wl[13221], wl[13222], wl[13223], wl[13224], wl[13225], wl[13226], wl[13227], wl[13228], wl[13229], wl[13230], wl[13231], wl[13232], wl[13233], wl[13234], wl[13235], wl[13236], wl[13237], wl[13238], wl[13239], wl[13240], wl[13241], wl[13242], wl[13243], wl[13244], wl[13245], wl[13246], wl[13247], wl[13248], wl[13249], wl[13250], wl[13251], wl[13252], wl[13253], wl[13254], wl[13255], wl[13256], wl[13257], wl[13258], wl[13259], wl[13260], wl[13261], wl[13262], wl[13263], wl[13264], wl[13265], wl[13266], wl[13267], wl[13268], wl[13269], wl[13270], wl[13271], wl[13272], wl[13273], wl[13274], wl[13275], wl[13276], wl[13277], wl[13278], wl[13279], wl[13280], wl[13281], wl[13282], wl[13283], wl[13284], wl[13285], wl[13286], wl[13287], wl[13288], wl[13289], wl[13290], wl[13291], wl[13292], wl[13293], wl[13294], wl[13295], wl[13296], wl[13297], wl[13298], wl[13299], wl[13300], wl[13301], wl[13302], wl[13303], wl[13304], wl[13305], wl[13306], wl[13307], wl[13308], wl[13309], wl[13310], wl[13311], wl[13312], wl[13313], wl[13314], wl[13315], wl[13316], wl[13317], wl[13318], wl[13319], wl[13320], wl[13321], wl[13322], wl[13323], wl[13324], wl[13325], wl[13326], wl[13327], wl[13328], wl[13329], wl[13330], wl[13331], wl[13332], wl[13333], wl[13334], wl[13335], wl[13336], wl[13337], wl[13338], wl[13339], wl[13340], wl[13341], wl[13342], wl[13343], wl[13344], wl[13345], wl[13346], wl[13347], wl[13348], wl[13349], wl[13350], wl[13351], wl[13352], wl[13353], wl[13354], wl[13355], wl[13356], wl[13357], wl[13358], wl[13359], wl[13360], wl[13361], wl[13362], wl[13363], wl[13364], wl[13365], wl[13366], wl[13367], wl[13368], wl[13369], wl[13370], wl[13371], wl[13372], wl[13373], wl[13374], wl[13375], wl[13376], wl[13377], wl[13378], wl[13379], wl[13380], wl[13381], wl[13382], wl[13383], wl[13384], wl[13385], wl[13386], wl[13387], wl[13388], wl[13389], wl[13390], wl[13391], wl[13392], wl[13393], wl[13394], wl[13395], wl[13396], wl[13397], wl[13398], wl[13399], wl[13400], wl[13401], wl[13402], wl[13403], wl[13404], wl[13405], wl[13406], wl[13407], wl[13408], wl[13409], wl[13410], wl[13411], wl[13412], wl[13413], wl[13414], wl[13415], wl[13416], wl[13417], wl[13418], wl[13419], wl[13420], wl[13421], wl[13422], wl[13423], wl[13424], wl[13425], wl[13426], wl[13427], wl[13428], wl[13429], wl[13430], wl[13431], wl[13432], wl[13433], wl[13434], wl[13435], wl[13436], wl[13437], wl[13438], wl[13439], wl[13440], wl[13441], wl[13442], wl[13443], wl[13444], wl[13445], wl[13446], wl[13447], wl[13448], wl[13449], wl[13450], wl[13451], wl[13452], wl[13453], wl[13454], wl[13455], wl[13456], wl[13457], wl[13458], wl[13459], wl[13460], wl[13461], wl[13462], wl[13463], wl[13464], wl[13465], wl[13466], wl[13467], wl[13468], wl[13469], wl[13470], wl[13471], wl[13472], wl[13473], wl[13474], wl[13475], wl[13476], wl[13477], wl[13478], wl[13479], wl[13480], wl[13481], wl[13482], wl[13483], wl[13484], wl[13485], wl[13486], wl[13487], wl[13488], wl[13489], wl[13490], wl[13491], wl[13492], wl[13493], wl[13494], wl[13495], wl[13496], wl[13497], wl[13498], wl[13499], wl[13500], wl[13501], wl[13502], wl[13503], wl[13504], wl[13505], wl[13506], wl[13507], wl[13508], wl[13509], wl[13510], wl[13511], wl[13512], wl[13513], wl[13514], wl[13515], wl[13516], wl[13517], wl[13518], wl[13519], wl[13520], wl[13521], wl[13522], wl[13523], wl[13524], wl[13525], wl[13526], wl[13527], wl[13528], wl[13529], wl[13530], wl[13531], wl[13532], wl[13533], wl[13534], wl[13535], wl[13536], wl[13537], wl[13538], wl[13539], wl[13540], wl[13541], wl[13542], wl[13543], wl[13544], wl[13545], wl[13546], wl[13547], wl[13548], wl[13549], wl[13550], wl[13551], wl[13552], wl[13553], wl[13554], wl[13555], wl[13556], wl[13557], wl[13558], wl[13559], wl[13560], wl[13561], wl[13562], wl[13563], wl[13564], wl[13565], wl[13566], wl[13567], wl[13568], wl[13569], wl[13570], wl[13571], wl[13572], wl[13573], wl[13574], wl[13575], wl[13576], wl[13577], wl[13578], wl[13579], wl[13580], wl[13581], wl[13582], wl[13583], wl[13584], wl[13585], wl[13586], wl[13587], wl[13588], wl[13589], wl[13590], wl[13591], wl[13592], wl[13593], wl[13594], wl[13595], wl[13596], wl[13597], wl[13598], wl[13599], wl[13600], wl[13601], wl[13602], wl[13603], wl[13604], wl[13605], wl[13606], wl[13607], wl[13608], wl[13609], wl[13610], wl[13611], wl[13612], wl[13613], wl[13614], wl[13615], wl[13616], wl[13617], wl[13618], wl[13619], wl[13620], wl[13621], wl[13622], wl[13623], wl[13624], wl[13625], wl[13626], wl[13627], wl[13628], wl[13629], wl[13630], wl[13631], wl[13632], wl[13633], wl[13634], wl[13635], wl[13636], wl[13637], wl[13638], wl[13639], wl[13640], wl[13641], wl[13642], wl[13643], wl[13644], wl[13645], wl[13646], wl[13647], wl[13648], wl[13649], wl[13650], wl[13651], wl[13652], wl[13653], wl[13654], wl[13655], wl[13656], wl[13657], wl[13658], wl[13659], wl[13660], wl[13661], wl[13662], wl[13663], wl[13664], wl[13665], wl[13666], wl[13667], wl[13668], wl[13669], wl[13670], wl[13671], wl[13672], wl[13673], wl[13674], wl[13675], wl[13676], wl[13677], wl[13678], wl[13679], wl[13680], wl[13681], wl[13682], wl[13683], wl[13684], wl[13685], wl[13686], wl[13687], wl[13688], wl[13689], wl[13690], wl[13691], wl[13692], wl[13693], wl[13694], wl[13695], wl[13696], wl[13697], wl[13698], wl[13699], wl[13700], wl[13701], wl[13702], wl[13703], wl[13704], wl[13705], wl[13706], wl[13707], wl[13708], wl[13709], wl[13710], wl[13711], wl[13712], wl[13713], wl[13714], wl[13715], wl[13716], wl[13717], wl[13718], wl[13719], wl[13720], wl[13721], wl[13722], wl[13723], wl[13724], wl[13725], wl[13726], wl[13727], wl[13728], wl[13729], wl[13730], wl[13731], wl[13732], wl[13733], wl[13734], wl[13735], wl[13736], wl[13737], wl[13738], wl[13739], wl[13740], wl[13741], wl[13742], wl[13743], wl[13744], wl[13745], wl[13746], wl[13747], wl[13748], wl[13749], wl[13750], wl[13751], wl[13752], wl[13753], wl[13754], wl[13755], wl[13756], wl[13757], wl[13758], wl[13759], wl[13760], wl[13761], wl[13762], wl[13763], wl[13764], wl[13765], wl[13766], wl[13767], wl[13768], wl[13769], wl[13770], wl[13771], wl[13772], wl[13773], wl[13774], wl[13775], wl[13776], wl[13777], wl[13778], wl[13779], wl[13780], wl[13781], wl[13782], wl[13783], wl[13784], wl[13785], wl[13786], wl[13787], wl[13788], wl[13789], wl[13790], wl[13791], wl[13792], wl[13793], wl[13794], wl[13795], wl[13796], wl[13797], wl[13798], wl[13799], wl[13800], wl[13801], wl[13802], wl[13803], wl[13804], wl[13805], wl[13806], wl[13807], wl[13808], wl[13809], wl[13810], wl[13811], wl[13812], wl[13813], wl[13814], wl[13815], wl[13816], wl[13817], wl[13818], wl[13819], wl[13820], wl[13821], wl[13822], wl[13823], wl[13824], wl[13825], wl[13826], wl[13827], wl[13828], wl[13829], wl[13830], wl[13831], wl[13832], wl[13833], wl[13834], wl[13835], wl[13836], wl[13837], wl[13838], wl[13839], wl[13840], wl[13841], wl[13842], wl[13843], wl[13844], wl[13845], wl[13846], wl[13847], wl[13848], wl[13849], wl[13850], wl[13851], wl[13852], wl[13853], wl[13854], wl[13855], wl[13856], wl[13857], wl[13858], wl[13859], wl[13860], wl[13861], wl[13862], wl[13863], wl[13864], wl[13865], wl[13866], wl[13867], wl[13868], wl[13869], wl[13870], wl[13871], wl[13872], wl[13873], wl[13874], wl[13875], wl[13876], wl[13877], wl[13878], wl[13879], wl[13880], wl[13881], wl[13882], wl[13883], wl[13884], wl[13885], wl[13886], wl[13887], wl[13888], wl[13889], wl[13890], wl[13891], wl[13892], wl[13893], wl[13894], wl[13895], wl[13896], wl[13897], wl[13898], wl[13899], wl[13900], wl[13901], wl[13902], wl[13903], wl[13904], wl[13905], wl[13906], wl[13907], wl[13908], wl[13909], wl[13910], wl[13911], wl[13912], wl[13913], wl[13914], wl[13915], wl[13916], wl[13917], wl[13918], wl[13919], wl[13920], wl[13921], wl[13922], wl[13923], wl[13924], wl[13925], wl[13926], wl[13927], wl[13928], wl[13929], wl[13930], wl[13931], wl[13932], wl[13933], wl[13934], wl[13935], wl[13936], wl[13937], wl[13938], wl[13939], wl[13940], wl[13941], wl[13942], wl[13943], wl[13944], wl[13945], wl[13946], wl[13947], wl[13948], wl[13949], wl[13950], wl[13951], wl[13952], wl[13953], wl[13954], wl[13955], wl[13956], wl[13957], wl[13958], wl[13959], wl[13960], wl[13961], wl[13962], wl[13963], wl[19068], wl[19069], wl[19070], wl[19071], wl[19072], wl[19073], wl[19074], wl[19075], wl[19076], wl[19077], wl[19078], wl[19079], wl[19080], wl[19081], wl[19082], wl[19083], wl[19084], wl[19085], wl[19086], wl[19087], wl[19088], wl[19089], wl[19090], wl[19091], wl[19092], wl[19093], wl[19094], wl[19095], wl[19096], wl[19097], wl[19098], wl[19099], wl[19100], wl[19101], wl[19102], wl[19103], wl[19104], wl[19105], wl[19106], wl[19107], wl[19108], wl[19109], wl[19110], wl[19111], wl[19112], wl[19113], wl[19114], wl[19115], wl[19116], wl[19117], wl[19118], wl[19119], wl[19120], wl[19121], wl[19122], wl[19123], wl[19124], wl[19125], wl[19126], wl[19127], wl[19128], wl[19129], wl[19130], wl[19131], wl[19132], wl[19133], wl[19134], wl[19135], wl[19136], wl[19137], wl[19138], wl[19139], wl[19140], wl[19141], wl[19142], wl[19143], wl[19144], wl[19145], wl[19146], wl[19147], wl[12864], wl[12865], wl[12866], wl[12867], wl[12868], wl[12869], wl[12870], wl[12871], wl[12872], wl[12873], wl[12874], wl[12875], wl[12876], wl[12877], wl[12878], wl[12879], wl[12880], wl[12881], wl[12882], wl[12883], wl[12884], wl[12885], wl[12886], wl[12887], wl[12888], wl[12889], wl[12890], wl[12891], wl[12892], wl[12893], wl[12894], wl[12895], wl[12896], wl[12897], wl[12898], wl[12899], wl[12900], wl[12901], wl[12902], wl[12903], wl[12904], wl[12905], wl[12906], wl[12907], wl[12908], wl[12909], wl[12910], wl[12911], wl[12912], wl[12913], wl[12914], wl[12915], wl[12916], wl[12917], wl[12918], wl[12919], wl[12920], wl[12921], wl[12922], wl[12923], wl[12924], wl[12925], wl[12926], wl[12927], wl[12928], wl[12929], wl[12930], wl[12931], wl[12932], wl[12933], wl[12934], wl[12935], wl[12936], wl[12937], wl[12938], wl[12939], wl[12940], wl[12941], wl[12942], wl[12943], wl[18988], wl[18989], wl[18990], wl[18991], wl[18992], wl[18993], wl[18994], wl[18995], wl[18996], wl[18997], wl[18998], wl[18999], wl[19000], wl[19001], wl[19002], wl[19003], wl[19004], wl[19005], wl[19006], wl[19007], wl[19008], wl[19009], wl[19010], wl[19011], wl[19012], wl[19013], wl[19014], wl[19015], wl[19016], wl[19017], wl[19018], wl[19019], wl[19020], wl[19021], wl[19022], wl[19023], wl[19024], wl[19025], wl[19026], wl[19027], wl[19028], wl[19029], wl[19030], wl[19031], wl[19032], wl[19033], wl[19034], wl[19035], wl[19036], wl[19037], wl[19038], wl[19039], wl[19040], wl[19041], wl[19042], wl[19043], wl[19044], wl[19045], wl[19046], wl[19047], wl[19048], wl[19049], wl[19050], wl[19051], wl[19052], wl[19053], wl[19054], wl[19055], wl[19056], wl[19057], wl[19058], wl[19059], wl[19060], wl[19061], wl[19062], wl[19063], wl[19064], wl[19065], wl[19066], wl[19067]})
    );
    tile tile_4__2_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_2__1__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_2__1__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_2__1__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_3__0__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_3__0__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_3__0__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_2__0__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_2__0__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_2__0__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_2__0__grid_top_r_in[1]),
        .grid_left_in(grid_clb_3__1__grid_left_in),
        .grid_bottom_in(grid_clb_3__1__grid_bottom_in),
        .chanx_left_in(sb_1__1__3_chanx_right_out),
        .chanx_left_out(cbx_1__1__6_chanx_left_out),
        .grid_top_out(grid_clb_3__2__grid_bottom_in),
        .chany_bottom_in(sb_1__0__2_chany_top_out),
        .chany_bottom_out(cby_1__1__8_chany_bottom_out),
        .grid_right_out(grid_clb_4__1__grid_left_in),
        .chany_top_in_0(cby_1__1__9_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__9_chanx_left_out),
        .chany_top_out_0(sb_1__1__6_chany_top_out),
        .chanx_right_out_0(sb_1__1__6_chanx_right_out),
        .grid_top_r_in(sb_3__1__grid_top_r_in),
        .grid_top_l_in(sb_3__1__grid_top_l_in),
        .grid_right_t_in(sb_3__1__grid_right_t_in),
        .grid_right_b_in(sb_3__1__grid_right_b_in),
        .grid_bottom_r_in(sb_3__0__grid_top_r_in),
        .grid_bottom_l_in(sb_3__0__grid_top_l_in),
        .grid_left_t_in(sb_2__1__grid_right_t_in),
        .grid_left_b_in(sb_2__1__grid_right_b_in),
        .bl({bl[4148], bl[4149], bl[4150], bl[4151], bl[4152], bl[4153], bl[4154], bl[4155], bl[4156], bl[4157], bl[4158], bl[4159], bl[4160], bl[4161], bl[4162], bl[4163], bl[4164], bl[4165], bl[4166], bl[4167], bl[4168], bl[4169], bl[4170], bl[4171], bl[4172], bl[4173], bl[4174], bl[4175], bl[4176], bl[4177], bl[4178], bl[4179], bl[4180], bl[4181], bl[4182], bl[4183], bl[4184], bl[4185], bl[4186], bl[4187], bl[4188], bl[4189], bl[4190], bl[4191], bl[4192], bl[4193], bl[4194], bl[4195], bl[4196], bl[4197], bl[4198], bl[4199], bl[4200], bl[4201], bl[4202], bl[4203], bl[4204], bl[4205], bl[4206], bl[4207], bl[4208], bl[4209], bl[4210], bl[4211], bl[4212], bl[4213], bl[4214], bl[4215], bl[4216], bl[4217], bl[4218], bl[4219], bl[4220], bl[4221], bl[4222], bl[4223], bl[4224], bl[4225], bl[4226], bl[4227], bl[4228], bl[4229], bl[4230], bl[4231], bl[4232], bl[4233], bl[4234], bl[4235], bl[4236], bl[4237], bl[4238], bl[4239], bl[4240], bl[4241], bl[4242], bl[4243], bl[4244], bl[4245], bl[4246], bl[4247], bl[4248], bl[4249], bl[4250], bl[4251], bl[4252], bl[4253], bl[4254], bl[4255], bl[4256], bl[4257], bl[4258], bl[4259], bl[4260], bl[4261], bl[4262], bl[4263], bl[4264], bl[4265], bl[4266], bl[4267], bl[4268], bl[4269], bl[4270], bl[4271], bl[4272], bl[4273], bl[4274], bl[4275], bl[4276], bl[4277], bl[4278], bl[4279], bl[4280], bl[4281], bl[4282], bl[4283], bl[4284], bl[4285], bl[4286], bl[4287], bl[4288], bl[4289], bl[4290], bl[4291], bl[4292], bl[4293], bl[4294], bl[4295], bl[4296], bl[4297], bl[4298], bl[4299], bl[4300], bl[4301], bl[4302], bl[4303], bl[4304], bl[4305], bl[4306], bl[4307], bl[4308], bl[4309], bl[4310], bl[4311], bl[4312], bl[4313], bl[4314], bl[4315], bl[4316], bl[4317], bl[4318], bl[4319], bl[4320], bl[4321], bl[4322], bl[4323], bl[4324], bl[4325], bl[4326], bl[4327], bl[4328], bl[4329], bl[4330], bl[4331], bl[4332], bl[4333], bl[4334], bl[4335], bl[4336], bl[4337], bl[4338], bl[4339], bl[4340], bl[4341], bl[4342], bl[4343], bl[4344], bl[4345], bl[4346], bl[4347], bl[4348], bl[4349], bl[4350], bl[4351], bl[4352], bl[4353], bl[4354], bl[4355], bl[4356], bl[4357], bl[4358], bl[4359], bl[4360], bl[4361], bl[4362], bl[4363], bl[4364], bl[4365], bl[4366], bl[4367], bl[4368], bl[4369], bl[4370], bl[4371], bl[4372], bl[4373], bl[4374], bl[4375], bl[4376], bl[4377], bl[4378], bl[4379], bl[4380], bl[4381], bl[4382], bl[4383], bl[4384], bl[4385], bl[4386], bl[4387], bl[4388], bl[4389], bl[4390], bl[4391], bl[4392], bl[4393], bl[4394], bl[4395], bl[4396], bl[4397], bl[4398], bl[4399], bl[4400], bl[4401], bl[4402], bl[4403], bl[4404], bl[4405], bl[4406], bl[4407], bl[4408], bl[4409], bl[4410], bl[4411], bl[4412], bl[4413], bl[4414], bl[4415], bl[4416], bl[4417], bl[4418], bl[4419], bl[4420], bl[4421], bl[4422], bl[4423], bl[4424], bl[4425], bl[4426], bl[4427], bl[4428], bl[4429], bl[4430], bl[4431], bl[4432], bl[4433], bl[4434], bl[4435], bl[4436], bl[4437], bl[4438], bl[4439], bl[4440], bl[4441], bl[4442], bl[4443], bl[4444], bl[4445], bl[4446], bl[4447], bl[4448], bl[4449], bl[4450], bl[4451], bl[4452], bl[4453], bl[4454], bl[4455], bl[4456], bl[4457], bl[4458], bl[4459], bl[4460], bl[4461], bl[4462], bl[4463], bl[4464], bl[4465], bl[4466], bl[4467], bl[4468], bl[4469], bl[4470], bl[4471], bl[4472], bl[4473], bl[4474], bl[4475], bl[4476], bl[4477], bl[4478], bl[4479], bl[4480], bl[4481], bl[4482], bl[4483], bl[4484], bl[4485], bl[4486], bl[4487], bl[4488], bl[4489], bl[4490], bl[4491], bl[4492], bl[4493], bl[4494], bl[4495], bl[4496], bl[4497], bl[4498], bl[4499], bl[4500], bl[4501], bl[4502], bl[4503], bl[4504], bl[4505], bl[4506], bl[4507], bl[4508], bl[4509], bl[4510], bl[4511], bl[4512], bl[4513], bl[4514], bl[4515], bl[4516], bl[4517], bl[4518], bl[4519], bl[4520], bl[4521], bl[4522], bl[4523], bl[4524], bl[4525], bl[4526], bl[4527], bl[4528], bl[4529], bl[4530], bl[4531], bl[4532], bl[4533], bl[4534], bl[4535], bl[4536], bl[4537], bl[4538], bl[4539], bl[4540], bl[4541], bl[4542], bl[4543], bl[4544], bl[4545], bl[4546], bl[4547], bl[4548], bl[4549], bl[4550], bl[4551], bl[4552], bl[4553], bl[4554], bl[4555], bl[4556], bl[4557], bl[4558], bl[4559], bl[4560], bl[4561], bl[4562], bl[4563], bl[4564], bl[4565], bl[4566], bl[4567], bl[4568], bl[4569], bl[4570], bl[4571], bl[4572], bl[4573], bl[4574], bl[4575], bl[4576], bl[4577], bl[4578], bl[4579], bl[4580], bl[4581], bl[4582], bl[4583], bl[4584], bl[4585], bl[4586], bl[4587], bl[4588], bl[4589], bl[4590], bl[4591], bl[4592], bl[4593], bl[4594], bl[4595], bl[4596], bl[4597], bl[4598], bl[4599], bl[4600], bl[4601], bl[4602], bl[4603], bl[4604], bl[4605], bl[4606], bl[4607], bl[4608], bl[4609], bl[4610], bl[4611], bl[4612], bl[4613], bl[4614], bl[4615], bl[4616], bl[4617], bl[4618], bl[4619], bl[4620], bl[4621], bl[4622], bl[4623], bl[4624], bl[4625], bl[4626], bl[4627], bl[4628], bl[4629], bl[4630], bl[4631], bl[4632], bl[4633], bl[4634], bl[4635], bl[4636], bl[4637], bl[4638], bl[4639], bl[4640], bl[4641], bl[4642], bl[4643], bl[4644], bl[4645], bl[4646], bl[4647], bl[4648], bl[4649], bl[4650], bl[4651], bl[4652], bl[4653], bl[4654], bl[4655], bl[4656], bl[4657], bl[4658], bl[4659], bl[4660], bl[4661], bl[4662], bl[4663], bl[4664], bl[4665], bl[4666], bl[4667], bl[4668], bl[4669], bl[4670], bl[4671], bl[4672], bl[4673], bl[4674], bl[4675], bl[4676], bl[4677], bl[4678], bl[4679], bl[4680], bl[4681], bl[4682], bl[4683], bl[4684], bl[4685], bl[4686], bl[4687], bl[4688], bl[4689], bl[4690], bl[4691], bl[4692], bl[4693], bl[4694], bl[4695], bl[4696], bl[4697], bl[4698], bl[4699], bl[4700], bl[4701], bl[4702], bl[4703], bl[4704], bl[4705], bl[4706], bl[4707], bl[4708], bl[4709], bl[4710], bl[4711], bl[4712], bl[4713], bl[4714], bl[4715], bl[4716], bl[4717], bl[4718], bl[4719], bl[4720], bl[4721], bl[4722], bl[4723], bl[4724], bl[4725], bl[4726], bl[4727], bl[4728], bl[4729], bl[4730], bl[4731], bl[4732], bl[4733], bl[4734], bl[4735], bl[4736], bl[4737], bl[4738], bl[4739], bl[4740], bl[4741], bl[4742], bl[4743], bl[4744], bl[4745], bl[4746], bl[4747], bl[4748], bl[4749], bl[4750], bl[4751], bl[4752], bl[4753], bl[4754], bl[4755], bl[4756], bl[4757], bl[4758], bl[4759], bl[4760], bl[4761], bl[4762], bl[4763], bl[4764], bl[4765], bl[4766], bl[4767], bl[4768], bl[4769], bl[4770], bl[4771], bl[4772], bl[4773], bl[4774], bl[4775], bl[4776], bl[4777], bl[4778], bl[4779], bl[4780], bl[4781], bl[4782], bl[4783], bl[4784], bl[4785], bl[4786], bl[4787], bl[4788], bl[4789], bl[4790], bl[4791], bl[4792], bl[4793], bl[4794], bl[4795], bl[4796], bl[4797], bl[4798], bl[4799], bl[4800], bl[4801], bl[4802], bl[4803], bl[4804], bl[4805], bl[4806], bl[4807], bl[4808], bl[4809], bl[4810], bl[4811], bl[4812], bl[4813], bl[4814], bl[4815], bl[4816], bl[4817], bl[4818], bl[4819], bl[4820], bl[4821], bl[4822], bl[4823], bl[4824], bl[4825], bl[4826], bl[4827], bl[4828], bl[4829], bl[4830], bl[4831], bl[4832], bl[4833], bl[4834], bl[4835], bl[4836], bl[4837], bl[4838], bl[4839], bl[4840], bl[4841], bl[4842], bl[4843], bl[4844], bl[4845], bl[4846], bl[4847], bl[4848], bl[4849], bl[4850], bl[4851], bl[4852], bl[4853], bl[4854], bl[4855], bl[4856], bl[4857], bl[4858], bl[4859], bl[4860], bl[4861], bl[4862], bl[4863], bl[4864], bl[4865], bl[4866], bl[4867], bl[4868], bl[4869], bl[4870], bl[4871], bl[4872], bl[4873], bl[4874], bl[4875], bl[4876], bl[4877], bl[4878], bl[4879], bl[4880], bl[4881], bl[4882], bl[4883], bl[4884], bl[4885], bl[4886], bl[4887], bl[4888], bl[4889], bl[4890], bl[4891], bl[4892], bl[4893], bl[4894], bl[4895], bl[4896], bl[4897], bl[4898], bl[4899], bl[4900], bl[4901], bl[4902], bl[4903], bl[4904], bl[4905], bl[4906], bl[4907], bl[4908], bl[4909], bl[4910], bl[4911], bl[4912], bl[4913], bl[4914], bl[4915], bl[4916], bl[4917], bl[4918], bl[4919], bl[4920], bl[4921], bl[4922], bl[4923], bl[4924], bl[4925], bl[4926], bl[4927], bl[4928], bl[4929], bl[4930], bl[4931], bl[4932], bl[4933], bl[4934], bl[4935], bl[4936], bl[4937], bl[4938], bl[4939], bl[4940], bl[4941], bl[4942], bl[4943], bl[4944], bl[4945], bl[4946], bl[4947], bl[4948], bl[4949], bl[4950], bl[4951], bl[4952], bl[4953], bl[4954], bl[4955], bl[4956], bl[4957], bl[4958], bl[4959], bl[4960], bl[4961], bl[4962], bl[4963], bl[4964], bl[4965], bl[4966], bl[4967], bl[4968], bl[4969], bl[4970], bl[4971], bl[4972], bl[4973], bl[4974], bl[4975], bl[4976], bl[4977], bl[4978], bl[4979], bl[4980], bl[4981], bl[4982], bl[4983], bl[4984], bl[4985], bl[4986], bl[4987], bl[4988], bl[4989], bl[4990], bl[4991], bl[4992], bl[4993], bl[4994], bl[4995], bl[4996], bl[4997], bl[4998], bl[4999], bl[5000], bl[5001], bl[5002], bl[5003], bl[5004], bl[5005], bl[5006], bl[5007], bl[5008], bl[5009], bl[5010], bl[5011], bl[5012], bl[5013], bl[5014], bl[5015], bl[5016], bl[5017], bl[5018], bl[5019], bl[5020], bl[5021], bl[5022], bl[5023], bl[5024], bl[5025], bl[5026], bl[5027], bl[5028], bl[5029], bl[5030], bl[5031], bl[5032], bl[5033], bl[5034], bl[5035], bl[5036], bl[5037], bl[5038], bl[5039], bl[5040], bl[5041], bl[5042], bl[5043], bl[5044], bl[5045], bl[5046], bl[5047], bl[5048], bl[5049], bl[5050], bl[5051], bl[5052], bl[5053], bl[5054], bl[5055], bl[5056], bl[5057], bl[5058], bl[5059], bl[5060], bl[5061], bl[5062], bl[5063], bl[5064], bl[5065], bl[5066], bl[5067], bl[5068], bl[5069], bl[5070], bl[5071], bl[5072], bl[5073], bl[5074], bl[5075], bl[5076], bl[5077], bl[5078], bl[5079], bl[5080], bl[5081], bl[5082], bl[5083], bl[5084], bl[5085], bl[5086], bl[5087], bl[5088], bl[5089], bl[5090], bl[5091], bl[5092], bl[5093], bl[5094], bl[5095], bl[5096], bl[5097], bl[5098], bl[5099], bl[5100], bl[5101], bl[5102], bl[5103], bl[5104], bl[5105], bl[5106], bl[5107], bl[5108], bl[5109], bl[5110], bl[5111], bl[5112], bl[5113], bl[5114], bl[5115], bl[5116], bl[5117], bl[5118], bl[5119], bl[5120], bl[5121], bl[5122], bl[5123], bl[5124], bl[5125], bl[5126], bl[5127], bl[5128], bl[5129], bl[5130], bl[5131], bl[5132], bl[5133], bl[5134], bl[5135], bl[5136], bl[5137], bl[5138], bl[5139], bl[5140], bl[5141], bl[5142], bl[5143], bl[5144], bl[5145], bl[5146], bl[5147], bl[5148], bl[5149], bl[5150], bl[5151], bl[5152], bl[5153], bl[5154], bl[5155], bl[5156], bl[5157], bl[5158], bl[5159], bl[5160], bl[5161], bl[5162], bl[5163], bl[5164], bl[5165], bl[5166], bl[5167], bl[7744], bl[7745], bl[7746], bl[7747], bl[7748], bl[7749], bl[7750], bl[7751], bl[7752], bl[7753], bl[7754], bl[7755], bl[7756], bl[7757], bl[7758], bl[7759], bl[7760], bl[7761], bl[7762], bl[7763], bl[7764], bl[7765], bl[7766], bl[7767], bl[7768], bl[7769], bl[7770], bl[7771], bl[7772], bl[7773], bl[7774], bl[7775], bl[7776], bl[7777], bl[7778], bl[7779], bl[7780], bl[7781], bl[7782], bl[7783], bl[7784], bl[7785], bl[7786], bl[7787], bl[7788], bl[7789], bl[7790], bl[7791], bl[7792], bl[7793], bl[7794], bl[7795], bl[7796], bl[7797], bl[7798], bl[7799], bl[7800], bl[7801], bl[7802], bl[7803], bl[7804], bl[7805], bl[7806], bl[7807], bl[7808], bl[7809], bl[7810], bl[7811], bl[7812], bl[7813], bl[7814], bl[7815], bl[7816], bl[7817], bl[7818], bl[7819], bl[7820], bl[7821], bl[7822], bl[7823], bl[4068], bl[4069], bl[4070], bl[4071], bl[4072], bl[4073], bl[4074], bl[4075], bl[4076], bl[4077], bl[4078], bl[4079], bl[4080], bl[4081], bl[4082], bl[4083], bl[4084], bl[4085], bl[4086], bl[4087], bl[4088], bl[4089], bl[4090], bl[4091], bl[4092], bl[4093], bl[4094], bl[4095], bl[4096], bl[4097], bl[4098], bl[4099], bl[4100], bl[4101], bl[4102], bl[4103], bl[4104], bl[4105], bl[4106], bl[4107], bl[4108], bl[4109], bl[4110], bl[4111], bl[4112], bl[4113], bl[4114], bl[4115], bl[4116], bl[4117], bl[4118], bl[4119], bl[4120], bl[4121], bl[4122], bl[4123], bl[4124], bl[4125], bl[4126], bl[4127], bl[4128], bl[4129], bl[4130], bl[4131], bl[4132], bl[4133], bl[4134], bl[4135], bl[4136], bl[4137], bl[4138], bl[4139], bl[4140], bl[4141], bl[4142], bl[4143], bl[4144], bl[4145], bl[4146], bl[4147], bl[7664], bl[7665], bl[7666], bl[7667], bl[7668], bl[7669], bl[7670], bl[7671], bl[7672], bl[7673], bl[7674], bl[7675], bl[7676], bl[7677], bl[7678], bl[7679], bl[7680], bl[7681], bl[7682], bl[7683], bl[7684], bl[7685], bl[7686], bl[7687], bl[7688], bl[7689], bl[7690], bl[7691], bl[7692], bl[7693], bl[7694], bl[7695], bl[7696], bl[7697], bl[7698], bl[7699], bl[7700], bl[7701], bl[7702], bl[7703], bl[7704], bl[7705], bl[7706], bl[7707], bl[7708], bl[7709], bl[7710], bl[7711], bl[7712], bl[7713], bl[7714], bl[7715], bl[7716], bl[7717], bl[7718], bl[7719], bl[7720], bl[7721], bl[7722], bl[7723], bl[7724], bl[7725], bl[7726], bl[7727], bl[7728], bl[7729], bl[7730], bl[7731], bl[7732], bl[7733], bl[7734], bl[7735], bl[7736], bl[7737], bl[7738], bl[7739], bl[7740], bl[7741], bl[7742], bl[7743]}),
        .wl({wl[4148], wl[4149], wl[4150], wl[4151], wl[4152], wl[4153], wl[4154], wl[4155], wl[4156], wl[4157], wl[4158], wl[4159], wl[4160], wl[4161], wl[4162], wl[4163], wl[4164], wl[4165], wl[4166], wl[4167], wl[4168], wl[4169], wl[4170], wl[4171], wl[4172], wl[4173], wl[4174], wl[4175], wl[4176], wl[4177], wl[4178], wl[4179], wl[4180], wl[4181], wl[4182], wl[4183], wl[4184], wl[4185], wl[4186], wl[4187], wl[4188], wl[4189], wl[4190], wl[4191], wl[4192], wl[4193], wl[4194], wl[4195], wl[4196], wl[4197], wl[4198], wl[4199], wl[4200], wl[4201], wl[4202], wl[4203], wl[4204], wl[4205], wl[4206], wl[4207], wl[4208], wl[4209], wl[4210], wl[4211], wl[4212], wl[4213], wl[4214], wl[4215], wl[4216], wl[4217], wl[4218], wl[4219], wl[4220], wl[4221], wl[4222], wl[4223], wl[4224], wl[4225], wl[4226], wl[4227], wl[4228], wl[4229], wl[4230], wl[4231], wl[4232], wl[4233], wl[4234], wl[4235], wl[4236], wl[4237], wl[4238], wl[4239], wl[4240], wl[4241], wl[4242], wl[4243], wl[4244], wl[4245], wl[4246], wl[4247], wl[4248], wl[4249], wl[4250], wl[4251], wl[4252], wl[4253], wl[4254], wl[4255], wl[4256], wl[4257], wl[4258], wl[4259], wl[4260], wl[4261], wl[4262], wl[4263], wl[4264], wl[4265], wl[4266], wl[4267], wl[4268], wl[4269], wl[4270], wl[4271], wl[4272], wl[4273], wl[4274], wl[4275], wl[4276], wl[4277], wl[4278], wl[4279], wl[4280], wl[4281], wl[4282], wl[4283], wl[4284], wl[4285], wl[4286], wl[4287], wl[4288], wl[4289], wl[4290], wl[4291], wl[4292], wl[4293], wl[4294], wl[4295], wl[4296], wl[4297], wl[4298], wl[4299], wl[4300], wl[4301], wl[4302], wl[4303], wl[4304], wl[4305], wl[4306], wl[4307], wl[4308], wl[4309], wl[4310], wl[4311], wl[4312], wl[4313], wl[4314], wl[4315], wl[4316], wl[4317], wl[4318], wl[4319], wl[4320], wl[4321], wl[4322], wl[4323], wl[4324], wl[4325], wl[4326], wl[4327], wl[4328], wl[4329], wl[4330], wl[4331], wl[4332], wl[4333], wl[4334], wl[4335], wl[4336], wl[4337], wl[4338], wl[4339], wl[4340], wl[4341], wl[4342], wl[4343], wl[4344], wl[4345], wl[4346], wl[4347], wl[4348], wl[4349], wl[4350], wl[4351], wl[4352], wl[4353], wl[4354], wl[4355], wl[4356], wl[4357], wl[4358], wl[4359], wl[4360], wl[4361], wl[4362], wl[4363], wl[4364], wl[4365], wl[4366], wl[4367], wl[4368], wl[4369], wl[4370], wl[4371], wl[4372], wl[4373], wl[4374], wl[4375], wl[4376], wl[4377], wl[4378], wl[4379], wl[4380], wl[4381], wl[4382], wl[4383], wl[4384], wl[4385], wl[4386], wl[4387], wl[4388], wl[4389], wl[4390], wl[4391], wl[4392], wl[4393], wl[4394], wl[4395], wl[4396], wl[4397], wl[4398], wl[4399], wl[4400], wl[4401], wl[4402], wl[4403], wl[4404], wl[4405], wl[4406], wl[4407], wl[4408], wl[4409], wl[4410], wl[4411], wl[4412], wl[4413], wl[4414], wl[4415], wl[4416], wl[4417], wl[4418], wl[4419], wl[4420], wl[4421], wl[4422], wl[4423], wl[4424], wl[4425], wl[4426], wl[4427], wl[4428], wl[4429], wl[4430], wl[4431], wl[4432], wl[4433], wl[4434], wl[4435], wl[4436], wl[4437], wl[4438], wl[4439], wl[4440], wl[4441], wl[4442], wl[4443], wl[4444], wl[4445], wl[4446], wl[4447], wl[4448], wl[4449], wl[4450], wl[4451], wl[4452], wl[4453], wl[4454], wl[4455], wl[4456], wl[4457], wl[4458], wl[4459], wl[4460], wl[4461], wl[4462], wl[4463], wl[4464], wl[4465], wl[4466], wl[4467], wl[4468], wl[4469], wl[4470], wl[4471], wl[4472], wl[4473], wl[4474], wl[4475], wl[4476], wl[4477], wl[4478], wl[4479], wl[4480], wl[4481], wl[4482], wl[4483], wl[4484], wl[4485], wl[4486], wl[4487], wl[4488], wl[4489], wl[4490], wl[4491], wl[4492], wl[4493], wl[4494], wl[4495], wl[4496], wl[4497], wl[4498], wl[4499], wl[4500], wl[4501], wl[4502], wl[4503], wl[4504], wl[4505], wl[4506], wl[4507], wl[4508], wl[4509], wl[4510], wl[4511], wl[4512], wl[4513], wl[4514], wl[4515], wl[4516], wl[4517], wl[4518], wl[4519], wl[4520], wl[4521], wl[4522], wl[4523], wl[4524], wl[4525], wl[4526], wl[4527], wl[4528], wl[4529], wl[4530], wl[4531], wl[4532], wl[4533], wl[4534], wl[4535], wl[4536], wl[4537], wl[4538], wl[4539], wl[4540], wl[4541], wl[4542], wl[4543], wl[4544], wl[4545], wl[4546], wl[4547], wl[4548], wl[4549], wl[4550], wl[4551], wl[4552], wl[4553], wl[4554], wl[4555], wl[4556], wl[4557], wl[4558], wl[4559], wl[4560], wl[4561], wl[4562], wl[4563], wl[4564], wl[4565], wl[4566], wl[4567], wl[4568], wl[4569], wl[4570], wl[4571], wl[4572], wl[4573], wl[4574], wl[4575], wl[4576], wl[4577], wl[4578], wl[4579], wl[4580], wl[4581], wl[4582], wl[4583], wl[4584], wl[4585], wl[4586], wl[4587], wl[4588], wl[4589], wl[4590], wl[4591], wl[4592], wl[4593], wl[4594], wl[4595], wl[4596], wl[4597], wl[4598], wl[4599], wl[4600], wl[4601], wl[4602], wl[4603], wl[4604], wl[4605], wl[4606], wl[4607], wl[4608], wl[4609], wl[4610], wl[4611], wl[4612], wl[4613], wl[4614], wl[4615], wl[4616], wl[4617], wl[4618], wl[4619], wl[4620], wl[4621], wl[4622], wl[4623], wl[4624], wl[4625], wl[4626], wl[4627], wl[4628], wl[4629], wl[4630], wl[4631], wl[4632], wl[4633], wl[4634], wl[4635], wl[4636], wl[4637], wl[4638], wl[4639], wl[4640], wl[4641], wl[4642], wl[4643], wl[4644], wl[4645], wl[4646], wl[4647], wl[4648], wl[4649], wl[4650], wl[4651], wl[4652], wl[4653], wl[4654], wl[4655], wl[4656], wl[4657], wl[4658], wl[4659], wl[4660], wl[4661], wl[4662], wl[4663], wl[4664], wl[4665], wl[4666], wl[4667], wl[4668], wl[4669], wl[4670], wl[4671], wl[4672], wl[4673], wl[4674], wl[4675], wl[4676], wl[4677], wl[4678], wl[4679], wl[4680], wl[4681], wl[4682], wl[4683], wl[4684], wl[4685], wl[4686], wl[4687], wl[4688], wl[4689], wl[4690], wl[4691], wl[4692], wl[4693], wl[4694], wl[4695], wl[4696], wl[4697], wl[4698], wl[4699], wl[4700], wl[4701], wl[4702], wl[4703], wl[4704], wl[4705], wl[4706], wl[4707], wl[4708], wl[4709], wl[4710], wl[4711], wl[4712], wl[4713], wl[4714], wl[4715], wl[4716], wl[4717], wl[4718], wl[4719], wl[4720], wl[4721], wl[4722], wl[4723], wl[4724], wl[4725], wl[4726], wl[4727], wl[4728], wl[4729], wl[4730], wl[4731], wl[4732], wl[4733], wl[4734], wl[4735], wl[4736], wl[4737], wl[4738], wl[4739], wl[4740], wl[4741], wl[4742], wl[4743], wl[4744], wl[4745], wl[4746], wl[4747], wl[4748], wl[4749], wl[4750], wl[4751], wl[4752], wl[4753], wl[4754], wl[4755], wl[4756], wl[4757], wl[4758], wl[4759], wl[4760], wl[4761], wl[4762], wl[4763], wl[4764], wl[4765], wl[4766], wl[4767], wl[4768], wl[4769], wl[4770], wl[4771], wl[4772], wl[4773], wl[4774], wl[4775], wl[4776], wl[4777], wl[4778], wl[4779], wl[4780], wl[4781], wl[4782], wl[4783], wl[4784], wl[4785], wl[4786], wl[4787], wl[4788], wl[4789], wl[4790], wl[4791], wl[4792], wl[4793], wl[4794], wl[4795], wl[4796], wl[4797], wl[4798], wl[4799], wl[4800], wl[4801], wl[4802], wl[4803], wl[4804], wl[4805], wl[4806], wl[4807], wl[4808], wl[4809], wl[4810], wl[4811], wl[4812], wl[4813], wl[4814], wl[4815], wl[4816], wl[4817], wl[4818], wl[4819], wl[4820], wl[4821], wl[4822], wl[4823], wl[4824], wl[4825], wl[4826], wl[4827], wl[4828], wl[4829], wl[4830], wl[4831], wl[4832], wl[4833], wl[4834], wl[4835], wl[4836], wl[4837], wl[4838], wl[4839], wl[4840], wl[4841], wl[4842], wl[4843], wl[4844], wl[4845], wl[4846], wl[4847], wl[4848], wl[4849], wl[4850], wl[4851], wl[4852], wl[4853], wl[4854], wl[4855], wl[4856], wl[4857], wl[4858], wl[4859], wl[4860], wl[4861], wl[4862], wl[4863], wl[4864], wl[4865], wl[4866], wl[4867], wl[4868], wl[4869], wl[4870], wl[4871], wl[4872], wl[4873], wl[4874], wl[4875], wl[4876], wl[4877], wl[4878], wl[4879], wl[4880], wl[4881], wl[4882], wl[4883], wl[4884], wl[4885], wl[4886], wl[4887], wl[4888], wl[4889], wl[4890], wl[4891], wl[4892], wl[4893], wl[4894], wl[4895], wl[4896], wl[4897], wl[4898], wl[4899], wl[4900], wl[4901], wl[4902], wl[4903], wl[4904], wl[4905], wl[4906], wl[4907], wl[4908], wl[4909], wl[4910], wl[4911], wl[4912], wl[4913], wl[4914], wl[4915], wl[4916], wl[4917], wl[4918], wl[4919], wl[4920], wl[4921], wl[4922], wl[4923], wl[4924], wl[4925], wl[4926], wl[4927], wl[4928], wl[4929], wl[4930], wl[4931], wl[4932], wl[4933], wl[4934], wl[4935], wl[4936], wl[4937], wl[4938], wl[4939], wl[4940], wl[4941], wl[4942], wl[4943], wl[4944], wl[4945], wl[4946], wl[4947], wl[4948], wl[4949], wl[4950], wl[4951], wl[4952], wl[4953], wl[4954], wl[4955], wl[4956], wl[4957], wl[4958], wl[4959], wl[4960], wl[4961], wl[4962], wl[4963], wl[4964], wl[4965], wl[4966], wl[4967], wl[4968], wl[4969], wl[4970], wl[4971], wl[4972], wl[4973], wl[4974], wl[4975], wl[4976], wl[4977], wl[4978], wl[4979], wl[4980], wl[4981], wl[4982], wl[4983], wl[4984], wl[4985], wl[4986], wl[4987], wl[4988], wl[4989], wl[4990], wl[4991], wl[4992], wl[4993], wl[4994], wl[4995], wl[4996], wl[4997], wl[4998], wl[4999], wl[5000], wl[5001], wl[5002], wl[5003], wl[5004], wl[5005], wl[5006], wl[5007], wl[5008], wl[5009], wl[5010], wl[5011], wl[5012], wl[5013], wl[5014], wl[5015], wl[5016], wl[5017], wl[5018], wl[5019], wl[5020], wl[5021], wl[5022], wl[5023], wl[5024], wl[5025], wl[5026], wl[5027], wl[5028], wl[5029], wl[5030], wl[5031], wl[5032], wl[5033], wl[5034], wl[5035], wl[5036], wl[5037], wl[5038], wl[5039], wl[5040], wl[5041], wl[5042], wl[5043], wl[5044], wl[5045], wl[5046], wl[5047], wl[5048], wl[5049], wl[5050], wl[5051], wl[5052], wl[5053], wl[5054], wl[5055], wl[5056], wl[5057], wl[5058], wl[5059], wl[5060], wl[5061], wl[5062], wl[5063], wl[5064], wl[5065], wl[5066], wl[5067], wl[5068], wl[5069], wl[5070], wl[5071], wl[5072], wl[5073], wl[5074], wl[5075], wl[5076], wl[5077], wl[5078], wl[5079], wl[5080], wl[5081], wl[5082], wl[5083], wl[5084], wl[5085], wl[5086], wl[5087], wl[5088], wl[5089], wl[5090], wl[5091], wl[5092], wl[5093], wl[5094], wl[5095], wl[5096], wl[5097], wl[5098], wl[5099], wl[5100], wl[5101], wl[5102], wl[5103], wl[5104], wl[5105], wl[5106], wl[5107], wl[5108], wl[5109], wl[5110], wl[5111], wl[5112], wl[5113], wl[5114], wl[5115], wl[5116], wl[5117], wl[5118], wl[5119], wl[5120], wl[5121], wl[5122], wl[5123], wl[5124], wl[5125], wl[5126], wl[5127], wl[5128], wl[5129], wl[5130], wl[5131], wl[5132], wl[5133], wl[5134], wl[5135], wl[5136], wl[5137], wl[5138], wl[5139], wl[5140], wl[5141], wl[5142], wl[5143], wl[5144], wl[5145], wl[5146], wl[5147], wl[5148], wl[5149], wl[5150], wl[5151], wl[5152], wl[5153], wl[5154], wl[5155], wl[5156], wl[5157], wl[5158], wl[5159], wl[5160], wl[5161], wl[5162], wl[5163], wl[5164], wl[5165], wl[5166], wl[5167], wl[7744], wl[7745], wl[7746], wl[7747], wl[7748], wl[7749], wl[7750], wl[7751], wl[7752], wl[7753], wl[7754], wl[7755], wl[7756], wl[7757], wl[7758], wl[7759], wl[7760], wl[7761], wl[7762], wl[7763], wl[7764], wl[7765], wl[7766], wl[7767], wl[7768], wl[7769], wl[7770], wl[7771], wl[7772], wl[7773], wl[7774], wl[7775], wl[7776], wl[7777], wl[7778], wl[7779], wl[7780], wl[7781], wl[7782], wl[7783], wl[7784], wl[7785], wl[7786], wl[7787], wl[7788], wl[7789], wl[7790], wl[7791], wl[7792], wl[7793], wl[7794], wl[7795], wl[7796], wl[7797], wl[7798], wl[7799], wl[7800], wl[7801], wl[7802], wl[7803], wl[7804], wl[7805], wl[7806], wl[7807], wl[7808], wl[7809], wl[7810], wl[7811], wl[7812], wl[7813], wl[7814], wl[7815], wl[7816], wl[7817], wl[7818], wl[7819], wl[7820], wl[7821], wl[7822], wl[7823], wl[4068], wl[4069], wl[4070], wl[4071], wl[4072], wl[4073], wl[4074], wl[4075], wl[4076], wl[4077], wl[4078], wl[4079], wl[4080], wl[4081], wl[4082], wl[4083], wl[4084], wl[4085], wl[4086], wl[4087], wl[4088], wl[4089], wl[4090], wl[4091], wl[4092], wl[4093], wl[4094], wl[4095], wl[4096], wl[4097], wl[4098], wl[4099], wl[4100], wl[4101], wl[4102], wl[4103], wl[4104], wl[4105], wl[4106], wl[4107], wl[4108], wl[4109], wl[4110], wl[4111], wl[4112], wl[4113], wl[4114], wl[4115], wl[4116], wl[4117], wl[4118], wl[4119], wl[4120], wl[4121], wl[4122], wl[4123], wl[4124], wl[4125], wl[4126], wl[4127], wl[4128], wl[4129], wl[4130], wl[4131], wl[4132], wl[4133], wl[4134], wl[4135], wl[4136], wl[4137], wl[4138], wl[4139], wl[4140], wl[4141], wl[4142], wl[4143], wl[4144], wl[4145], wl[4146], wl[4147], wl[7664], wl[7665], wl[7666], wl[7667], wl[7668], wl[7669], wl[7670], wl[7671], wl[7672], wl[7673], wl[7674], wl[7675], wl[7676], wl[7677], wl[7678], wl[7679], wl[7680], wl[7681], wl[7682], wl[7683], wl[7684], wl[7685], wl[7686], wl[7687], wl[7688], wl[7689], wl[7690], wl[7691], wl[7692], wl[7693], wl[7694], wl[7695], wl[7696], wl[7697], wl[7698], wl[7699], wl[7700], wl[7701], wl[7702], wl[7703], wl[7704], wl[7705], wl[7706], wl[7707], wl[7708], wl[7709], wl[7710], wl[7711], wl[7712], wl[7713], wl[7714], wl[7715], wl[7716], wl[7717], wl[7718], wl[7719], wl[7720], wl[7721], wl[7722], wl[7723], wl[7724], wl[7725], wl[7726], wl[7727], wl[7728], wl[7729], wl[7730], wl[7731], wl[7732], wl[7733], wl[7734], wl[7735], wl[7736], wl[7737], wl[7738], wl[7739], wl[7740], wl[7741], wl[7742], wl[7743]})
    );
    tile tile_4__3_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_2__2__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_2__2__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_2__2__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_3__1__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_3__1__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_3__1__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_2__1__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_2__1__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_2__1__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_2__1__grid_top_r_in[1]),
        .grid_left_in(grid_clb_3__2__grid_left_in),
        .grid_bottom_in(grid_clb_3__2__grid_bottom_in),
        .chanx_left_in(sb_1__1__4_chanx_right_out),
        .chanx_left_out(cbx_1__1__7_chanx_left_out),
        .grid_top_out(grid_clb_3__3__grid_bottom_in),
        .chany_bottom_in(sb_1__1__6_chany_top_out),
        .chany_bottom_out(cby_1__1__9_chany_bottom_out),
        .grid_right_out(grid_clb_4__2__grid_left_in),
        .chany_top_in_0(cby_1__1__10_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__10_chanx_left_out),
        .chany_top_out_0(sb_1__1__7_chany_top_out),
        .chanx_right_out_0(sb_1__1__7_chanx_right_out),
        .grid_top_r_in(sb_3__2__grid_top_r_in),
        .grid_top_l_in(sb_3__2__grid_top_l_in),
        .grid_right_t_in(sb_3__2__grid_right_t_in),
        .grid_right_b_in(sb_3__2__grid_right_b_in),
        .grid_bottom_r_in(sb_3__1__grid_top_r_in),
        .grid_bottom_l_in(sb_3__1__grid_top_l_in),
        .grid_left_t_in(sb_2__2__grid_right_t_in),
        .grid_left_b_in(sb_2__2__grid_right_b_in),
        .bl({bl[7904], bl[7905], bl[7906], bl[7907], bl[7908], bl[7909], bl[7910], bl[7911], bl[7912], bl[7913], bl[7914], bl[7915], bl[7916], bl[7917], bl[7918], bl[7919], bl[7920], bl[7921], bl[7922], bl[7923], bl[7924], bl[7925], bl[7926], bl[7927], bl[7928], bl[7929], bl[7930], bl[7931], bl[7932], bl[7933], bl[7934], bl[7935], bl[7936], bl[7937], bl[7938], bl[7939], bl[7940], bl[7941], bl[7942], bl[7943], bl[7944], bl[7945], bl[7946], bl[7947], bl[7948], bl[7949], bl[7950], bl[7951], bl[7952], bl[7953], bl[7954], bl[7955], bl[7956], bl[7957], bl[7958], bl[7959], bl[7960], bl[7961], bl[7962], bl[7963], bl[7964], bl[7965], bl[7966], bl[7967], bl[7968], bl[7969], bl[7970], bl[7971], bl[7972], bl[7973], bl[7974], bl[7975], bl[7976], bl[7977], bl[7978], bl[7979], bl[7980], bl[7981], bl[7982], bl[7983], bl[7984], bl[7985], bl[7986], bl[7987], bl[7988], bl[7989], bl[7990], bl[7991], bl[7992], bl[7993], bl[7994], bl[7995], bl[7996], bl[7997], bl[7998], bl[7999], bl[8000], bl[8001], bl[8002], bl[8003], bl[8004], bl[8005], bl[8006], bl[8007], bl[8008], bl[8009], bl[8010], bl[8011], bl[8012], bl[8013], bl[8014], bl[8015], bl[8016], bl[8017], bl[8018], bl[8019], bl[8020], bl[8021], bl[8022], bl[8023], bl[8024], bl[8025], bl[8026], bl[8027], bl[8028], bl[8029], bl[8030], bl[8031], bl[8032], bl[8033], bl[8034], bl[8035], bl[8036], bl[8037], bl[8038], bl[8039], bl[8040], bl[8041], bl[8042], bl[8043], bl[8044], bl[8045], bl[8046], bl[8047], bl[8048], bl[8049], bl[8050], bl[8051], bl[8052], bl[8053], bl[8054], bl[8055], bl[8056], bl[8057], bl[8058], bl[8059], bl[8060], bl[8061], bl[8062], bl[8063], bl[8064], bl[8065], bl[8066], bl[8067], bl[8068], bl[8069], bl[8070], bl[8071], bl[8072], bl[8073], bl[8074], bl[8075], bl[8076], bl[8077], bl[8078], bl[8079], bl[8080], bl[8081], bl[8082], bl[8083], bl[8084], bl[8085], bl[8086], bl[8087], bl[8088], bl[8089], bl[8090], bl[8091], bl[8092], bl[8093], bl[8094], bl[8095], bl[8096], bl[8097], bl[8098], bl[8099], bl[8100], bl[8101], bl[8102], bl[8103], bl[8104], bl[8105], bl[8106], bl[8107], bl[8108], bl[8109], bl[8110], bl[8111], bl[8112], bl[8113], bl[8114], bl[8115], bl[8116], bl[8117], bl[8118], bl[8119], bl[8120], bl[8121], bl[8122], bl[8123], bl[8124], bl[8125], bl[8126], bl[8127], bl[8128], bl[8129], bl[8130], bl[8131], bl[8132], bl[8133], bl[8134], bl[8135], bl[8136], bl[8137], bl[8138], bl[8139], bl[8140], bl[8141], bl[8142], bl[8143], bl[8144], bl[8145], bl[8146], bl[8147], bl[8148], bl[8149], bl[8150], bl[8151], bl[8152], bl[8153], bl[8154], bl[8155], bl[8156], bl[8157], bl[8158], bl[8159], bl[8160], bl[8161], bl[8162], bl[8163], bl[8164], bl[8165], bl[8166], bl[8167], bl[8168], bl[8169], bl[8170], bl[8171], bl[8172], bl[8173], bl[8174], bl[8175], bl[8176], bl[8177], bl[8178], bl[8179], bl[8180], bl[8181], bl[8182], bl[8183], bl[8184], bl[8185], bl[8186], bl[8187], bl[8188], bl[8189], bl[8190], bl[8191], bl[8192], bl[8193], bl[8194], bl[8195], bl[8196], bl[8197], bl[8198], bl[8199], bl[8200], bl[8201], bl[8202], bl[8203], bl[8204], bl[8205], bl[8206], bl[8207], bl[8208], bl[8209], bl[8210], bl[8211], bl[8212], bl[8213], bl[8214], bl[8215], bl[8216], bl[8217], bl[8218], bl[8219], bl[8220], bl[8221], bl[8222], bl[8223], bl[8224], bl[8225], bl[8226], bl[8227], bl[8228], bl[8229], bl[8230], bl[8231], bl[8232], bl[8233], bl[8234], bl[8235], bl[8236], bl[8237], bl[8238], bl[8239], bl[8240], bl[8241], bl[8242], bl[8243], bl[8244], bl[8245], bl[8246], bl[8247], bl[8248], bl[8249], bl[8250], bl[8251], bl[8252], bl[8253], bl[8254], bl[8255], bl[8256], bl[8257], bl[8258], bl[8259], bl[8260], bl[8261], bl[8262], bl[8263], bl[8264], bl[8265], bl[8266], bl[8267], bl[8268], bl[8269], bl[8270], bl[8271], bl[8272], bl[8273], bl[8274], bl[8275], bl[8276], bl[8277], bl[8278], bl[8279], bl[8280], bl[8281], bl[8282], bl[8283], bl[8284], bl[8285], bl[8286], bl[8287], bl[8288], bl[8289], bl[8290], bl[8291], bl[8292], bl[8293], bl[8294], bl[8295], bl[8296], bl[8297], bl[8298], bl[8299], bl[8300], bl[8301], bl[8302], bl[8303], bl[8304], bl[8305], bl[8306], bl[8307], bl[8308], bl[8309], bl[8310], bl[8311], bl[8312], bl[8313], bl[8314], bl[8315], bl[8316], bl[8317], bl[8318], bl[8319], bl[8320], bl[8321], bl[8322], bl[8323], bl[8324], bl[8325], bl[8326], bl[8327], bl[8328], bl[8329], bl[8330], bl[8331], bl[8332], bl[8333], bl[8334], bl[8335], bl[8336], bl[8337], bl[8338], bl[8339], bl[8340], bl[8341], bl[8342], bl[8343], bl[8344], bl[8345], bl[8346], bl[8347], bl[8348], bl[8349], bl[8350], bl[8351], bl[8352], bl[8353], bl[8354], bl[8355], bl[8356], bl[8357], bl[8358], bl[8359], bl[8360], bl[8361], bl[8362], bl[8363], bl[8364], bl[8365], bl[8366], bl[8367], bl[8368], bl[8369], bl[8370], bl[8371], bl[8372], bl[8373], bl[8374], bl[8375], bl[8376], bl[8377], bl[8378], bl[8379], bl[8380], bl[8381], bl[8382], bl[8383], bl[8384], bl[8385], bl[8386], bl[8387], bl[8388], bl[8389], bl[8390], bl[8391], bl[8392], bl[8393], bl[8394], bl[8395], bl[8396], bl[8397], bl[8398], bl[8399], bl[8400], bl[8401], bl[8402], bl[8403], bl[8404], bl[8405], bl[8406], bl[8407], bl[8408], bl[8409], bl[8410], bl[8411], bl[8412], bl[8413], bl[8414], bl[8415], bl[8416], bl[8417], bl[8418], bl[8419], bl[8420], bl[8421], bl[8422], bl[8423], bl[8424], bl[8425], bl[8426], bl[8427], bl[8428], bl[8429], bl[8430], bl[8431], bl[8432], bl[8433], bl[8434], bl[8435], bl[8436], bl[8437], bl[8438], bl[8439], bl[8440], bl[8441], bl[8442], bl[8443], bl[8444], bl[8445], bl[8446], bl[8447], bl[8448], bl[8449], bl[8450], bl[8451], bl[8452], bl[8453], bl[8454], bl[8455], bl[8456], bl[8457], bl[8458], bl[8459], bl[8460], bl[8461], bl[8462], bl[8463], bl[8464], bl[8465], bl[8466], bl[8467], bl[8468], bl[8469], bl[8470], bl[8471], bl[8472], bl[8473], bl[8474], bl[8475], bl[8476], bl[8477], bl[8478], bl[8479], bl[8480], bl[8481], bl[8482], bl[8483], bl[8484], bl[8485], bl[8486], bl[8487], bl[8488], bl[8489], bl[8490], bl[8491], bl[8492], bl[8493], bl[8494], bl[8495], bl[8496], bl[8497], bl[8498], bl[8499], bl[8500], bl[8501], bl[8502], bl[8503], bl[8504], bl[8505], bl[8506], bl[8507], bl[8508], bl[8509], bl[8510], bl[8511], bl[8512], bl[8513], bl[8514], bl[8515], bl[8516], bl[8517], bl[8518], bl[8519], bl[8520], bl[8521], bl[8522], bl[8523], bl[8524], bl[8525], bl[8526], bl[8527], bl[8528], bl[8529], bl[8530], bl[8531], bl[8532], bl[8533], bl[8534], bl[8535], bl[8536], bl[8537], bl[8538], bl[8539], bl[8540], bl[8541], bl[8542], bl[8543], bl[8544], bl[8545], bl[8546], bl[8547], bl[8548], bl[8549], bl[8550], bl[8551], bl[8552], bl[8553], bl[8554], bl[8555], bl[8556], bl[8557], bl[8558], bl[8559], bl[8560], bl[8561], bl[8562], bl[8563], bl[8564], bl[8565], bl[8566], bl[8567], bl[8568], bl[8569], bl[8570], bl[8571], bl[8572], bl[8573], bl[8574], bl[8575], bl[8576], bl[8577], bl[8578], bl[8579], bl[8580], bl[8581], bl[8582], bl[8583], bl[8584], bl[8585], bl[8586], bl[8587], bl[8588], bl[8589], bl[8590], bl[8591], bl[8592], bl[8593], bl[8594], bl[8595], bl[8596], bl[8597], bl[8598], bl[8599], bl[8600], bl[8601], bl[8602], bl[8603], bl[8604], bl[8605], bl[8606], bl[8607], bl[8608], bl[8609], bl[8610], bl[8611], bl[8612], bl[8613], bl[8614], bl[8615], bl[8616], bl[8617], bl[8618], bl[8619], bl[8620], bl[8621], bl[8622], bl[8623], bl[8624], bl[8625], bl[8626], bl[8627], bl[8628], bl[8629], bl[8630], bl[8631], bl[8632], bl[8633], bl[8634], bl[8635], bl[8636], bl[8637], bl[8638], bl[8639], bl[8640], bl[8641], bl[8642], bl[8643], bl[8644], bl[8645], bl[8646], bl[8647], bl[8648], bl[8649], bl[8650], bl[8651], bl[8652], bl[8653], bl[8654], bl[8655], bl[8656], bl[8657], bl[8658], bl[8659], bl[8660], bl[8661], bl[8662], bl[8663], bl[8664], bl[8665], bl[8666], bl[8667], bl[8668], bl[8669], bl[8670], bl[8671], bl[8672], bl[8673], bl[8674], bl[8675], bl[8676], bl[8677], bl[8678], bl[8679], bl[8680], bl[8681], bl[8682], bl[8683], bl[8684], bl[8685], bl[8686], bl[8687], bl[8688], bl[8689], bl[8690], bl[8691], bl[8692], bl[8693], bl[8694], bl[8695], bl[8696], bl[8697], bl[8698], bl[8699], bl[8700], bl[8701], bl[8702], bl[8703], bl[8704], bl[8705], bl[8706], bl[8707], bl[8708], bl[8709], bl[8710], bl[8711], bl[8712], bl[8713], bl[8714], bl[8715], bl[8716], bl[8717], bl[8718], bl[8719], bl[8720], bl[8721], bl[8722], bl[8723], bl[8724], bl[8725], bl[8726], bl[8727], bl[8728], bl[8729], bl[8730], bl[8731], bl[8732], bl[8733], bl[8734], bl[8735], bl[8736], bl[8737], bl[8738], bl[8739], bl[8740], bl[8741], bl[8742], bl[8743], bl[8744], bl[8745], bl[8746], bl[8747], bl[8748], bl[8749], bl[8750], bl[8751], bl[8752], bl[8753], bl[8754], bl[8755], bl[8756], bl[8757], bl[8758], bl[8759], bl[8760], bl[8761], bl[8762], bl[8763], bl[8764], bl[8765], bl[8766], bl[8767], bl[8768], bl[8769], bl[8770], bl[8771], bl[8772], bl[8773], bl[8774], bl[8775], bl[8776], bl[8777], bl[8778], bl[8779], bl[8780], bl[8781], bl[8782], bl[8783], bl[8784], bl[8785], bl[8786], bl[8787], bl[8788], bl[8789], bl[8790], bl[8791], bl[8792], bl[8793], bl[8794], bl[8795], bl[8796], bl[8797], bl[8798], bl[8799], bl[8800], bl[8801], bl[8802], bl[8803], bl[8804], bl[8805], bl[8806], bl[8807], bl[8808], bl[8809], bl[8810], bl[8811], bl[8812], bl[8813], bl[8814], bl[8815], bl[8816], bl[8817], bl[8818], bl[8819], bl[8820], bl[8821], bl[8822], bl[8823], bl[8824], bl[8825], bl[8826], bl[8827], bl[8828], bl[8829], bl[8830], bl[8831], bl[8832], bl[8833], bl[8834], bl[8835], bl[8836], bl[8837], bl[8838], bl[8839], bl[8840], bl[8841], bl[8842], bl[8843], bl[8844], bl[8845], bl[8846], bl[8847], bl[8848], bl[8849], bl[8850], bl[8851], bl[8852], bl[8853], bl[8854], bl[8855], bl[8856], bl[8857], bl[8858], bl[8859], bl[8860], bl[8861], bl[8862], bl[8863], bl[8864], bl[8865], bl[8866], bl[8867], bl[8868], bl[8869], bl[8870], bl[8871], bl[8872], bl[8873], bl[8874], bl[8875], bl[8876], bl[8877], bl[8878], bl[8879], bl[8880], bl[8881], bl[8882], bl[8883], bl[8884], bl[8885], bl[8886], bl[8887], bl[8888], bl[8889], bl[8890], bl[8891], bl[8892], bl[8893], bl[8894], bl[8895], bl[8896], bl[8897], bl[8898], bl[8899], bl[8900], bl[8901], bl[8902], bl[8903], bl[8904], bl[8905], bl[8906], bl[8907], bl[8908], bl[8909], bl[8910], bl[8911], bl[8912], bl[8913], bl[8914], bl[8915], bl[8916], bl[8917], bl[8918], bl[8919], bl[8920], bl[8921], bl[8922], bl[8923], bl[14044], bl[14045], bl[14046], bl[14047], bl[14048], bl[14049], bl[14050], bl[14051], bl[14052], bl[14053], bl[14054], bl[14055], bl[14056], bl[14057], bl[14058], bl[14059], bl[14060], bl[14061], bl[14062], bl[14063], bl[14064], bl[14065], bl[14066], bl[14067], bl[14068], bl[14069], bl[14070], bl[14071], bl[14072], bl[14073], bl[14074], bl[14075], bl[14076], bl[14077], bl[14078], bl[14079], bl[14080], bl[14081], bl[14082], bl[14083], bl[14084], bl[14085], bl[14086], bl[14087], bl[14088], bl[14089], bl[14090], bl[14091], bl[14092], bl[14093], bl[14094], bl[14095], bl[14096], bl[14097], bl[14098], bl[14099], bl[14100], bl[14101], bl[14102], bl[14103], bl[14104], bl[14105], bl[14106], bl[14107], bl[14108], bl[14109], bl[14110], bl[14111], bl[14112], bl[14113], bl[14114], bl[14115], bl[14116], bl[14117], bl[14118], bl[14119], bl[14120], bl[14121], bl[14122], bl[14123], bl[7824], bl[7825], bl[7826], bl[7827], bl[7828], bl[7829], bl[7830], bl[7831], bl[7832], bl[7833], bl[7834], bl[7835], bl[7836], bl[7837], bl[7838], bl[7839], bl[7840], bl[7841], bl[7842], bl[7843], bl[7844], bl[7845], bl[7846], bl[7847], bl[7848], bl[7849], bl[7850], bl[7851], bl[7852], bl[7853], bl[7854], bl[7855], bl[7856], bl[7857], bl[7858], bl[7859], bl[7860], bl[7861], bl[7862], bl[7863], bl[7864], bl[7865], bl[7866], bl[7867], bl[7868], bl[7869], bl[7870], bl[7871], bl[7872], bl[7873], bl[7874], bl[7875], bl[7876], bl[7877], bl[7878], bl[7879], bl[7880], bl[7881], bl[7882], bl[7883], bl[7884], bl[7885], bl[7886], bl[7887], bl[7888], bl[7889], bl[7890], bl[7891], bl[7892], bl[7893], bl[7894], bl[7895], bl[7896], bl[7897], bl[7898], bl[7899], bl[7900], bl[7901], bl[7902], bl[7903], bl[13964], bl[13965], bl[13966], bl[13967], bl[13968], bl[13969], bl[13970], bl[13971], bl[13972], bl[13973], bl[13974], bl[13975], bl[13976], bl[13977], bl[13978], bl[13979], bl[13980], bl[13981], bl[13982], bl[13983], bl[13984], bl[13985], bl[13986], bl[13987], bl[13988], bl[13989], bl[13990], bl[13991], bl[13992], bl[13993], bl[13994], bl[13995], bl[13996], bl[13997], bl[13998], bl[13999], bl[14000], bl[14001], bl[14002], bl[14003], bl[14004], bl[14005], bl[14006], bl[14007], bl[14008], bl[14009], bl[14010], bl[14011], bl[14012], bl[14013], bl[14014], bl[14015], bl[14016], bl[14017], bl[14018], bl[14019], bl[14020], bl[14021], bl[14022], bl[14023], bl[14024], bl[14025], bl[14026], bl[14027], bl[14028], bl[14029], bl[14030], bl[14031], bl[14032], bl[14033], bl[14034], bl[14035], bl[14036], bl[14037], bl[14038], bl[14039], bl[14040], bl[14041], bl[14042], bl[14043]}),
        .wl({wl[7904], wl[7905], wl[7906], wl[7907], wl[7908], wl[7909], wl[7910], wl[7911], wl[7912], wl[7913], wl[7914], wl[7915], wl[7916], wl[7917], wl[7918], wl[7919], wl[7920], wl[7921], wl[7922], wl[7923], wl[7924], wl[7925], wl[7926], wl[7927], wl[7928], wl[7929], wl[7930], wl[7931], wl[7932], wl[7933], wl[7934], wl[7935], wl[7936], wl[7937], wl[7938], wl[7939], wl[7940], wl[7941], wl[7942], wl[7943], wl[7944], wl[7945], wl[7946], wl[7947], wl[7948], wl[7949], wl[7950], wl[7951], wl[7952], wl[7953], wl[7954], wl[7955], wl[7956], wl[7957], wl[7958], wl[7959], wl[7960], wl[7961], wl[7962], wl[7963], wl[7964], wl[7965], wl[7966], wl[7967], wl[7968], wl[7969], wl[7970], wl[7971], wl[7972], wl[7973], wl[7974], wl[7975], wl[7976], wl[7977], wl[7978], wl[7979], wl[7980], wl[7981], wl[7982], wl[7983], wl[7984], wl[7985], wl[7986], wl[7987], wl[7988], wl[7989], wl[7990], wl[7991], wl[7992], wl[7993], wl[7994], wl[7995], wl[7996], wl[7997], wl[7998], wl[7999], wl[8000], wl[8001], wl[8002], wl[8003], wl[8004], wl[8005], wl[8006], wl[8007], wl[8008], wl[8009], wl[8010], wl[8011], wl[8012], wl[8013], wl[8014], wl[8015], wl[8016], wl[8017], wl[8018], wl[8019], wl[8020], wl[8021], wl[8022], wl[8023], wl[8024], wl[8025], wl[8026], wl[8027], wl[8028], wl[8029], wl[8030], wl[8031], wl[8032], wl[8033], wl[8034], wl[8035], wl[8036], wl[8037], wl[8038], wl[8039], wl[8040], wl[8041], wl[8042], wl[8043], wl[8044], wl[8045], wl[8046], wl[8047], wl[8048], wl[8049], wl[8050], wl[8051], wl[8052], wl[8053], wl[8054], wl[8055], wl[8056], wl[8057], wl[8058], wl[8059], wl[8060], wl[8061], wl[8062], wl[8063], wl[8064], wl[8065], wl[8066], wl[8067], wl[8068], wl[8069], wl[8070], wl[8071], wl[8072], wl[8073], wl[8074], wl[8075], wl[8076], wl[8077], wl[8078], wl[8079], wl[8080], wl[8081], wl[8082], wl[8083], wl[8084], wl[8085], wl[8086], wl[8087], wl[8088], wl[8089], wl[8090], wl[8091], wl[8092], wl[8093], wl[8094], wl[8095], wl[8096], wl[8097], wl[8098], wl[8099], wl[8100], wl[8101], wl[8102], wl[8103], wl[8104], wl[8105], wl[8106], wl[8107], wl[8108], wl[8109], wl[8110], wl[8111], wl[8112], wl[8113], wl[8114], wl[8115], wl[8116], wl[8117], wl[8118], wl[8119], wl[8120], wl[8121], wl[8122], wl[8123], wl[8124], wl[8125], wl[8126], wl[8127], wl[8128], wl[8129], wl[8130], wl[8131], wl[8132], wl[8133], wl[8134], wl[8135], wl[8136], wl[8137], wl[8138], wl[8139], wl[8140], wl[8141], wl[8142], wl[8143], wl[8144], wl[8145], wl[8146], wl[8147], wl[8148], wl[8149], wl[8150], wl[8151], wl[8152], wl[8153], wl[8154], wl[8155], wl[8156], wl[8157], wl[8158], wl[8159], wl[8160], wl[8161], wl[8162], wl[8163], wl[8164], wl[8165], wl[8166], wl[8167], wl[8168], wl[8169], wl[8170], wl[8171], wl[8172], wl[8173], wl[8174], wl[8175], wl[8176], wl[8177], wl[8178], wl[8179], wl[8180], wl[8181], wl[8182], wl[8183], wl[8184], wl[8185], wl[8186], wl[8187], wl[8188], wl[8189], wl[8190], wl[8191], wl[8192], wl[8193], wl[8194], wl[8195], wl[8196], wl[8197], wl[8198], wl[8199], wl[8200], wl[8201], wl[8202], wl[8203], wl[8204], wl[8205], wl[8206], wl[8207], wl[8208], wl[8209], wl[8210], wl[8211], wl[8212], wl[8213], wl[8214], wl[8215], wl[8216], wl[8217], wl[8218], wl[8219], wl[8220], wl[8221], wl[8222], wl[8223], wl[8224], wl[8225], wl[8226], wl[8227], wl[8228], wl[8229], wl[8230], wl[8231], wl[8232], wl[8233], wl[8234], wl[8235], wl[8236], wl[8237], wl[8238], wl[8239], wl[8240], wl[8241], wl[8242], wl[8243], wl[8244], wl[8245], wl[8246], wl[8247], wl[8248], wl[8249], wl[8250], wl[8251], wl[8252], wl[8253], wl[8254], wl[8255], wl[8256], wl[8257], wl[8258], wl[8259], wl[8260], wl[8261], wl[8262], wl[8263], wl[8264], wl[8265], wl[8266], wl[8267], wl[8268], wl[8269], wl[8270], wl[8271], wl[8272], wl[8273], wl[8274], wl[8275], wl[8276], wl[8277], wl[8278], wl[8279], wl[8280], wl[8281], wl[8282], wl[8283], wl[8284], wl[8285], wl[8286], wl[8287], wl[8288], wl[8289], wl[8290], wl[8291], wl[8292], wl[8293], wl[8294], wl[8295], wl[8296], wl[8297], wl[8298], wl[8299], wl[8300], wl[8301], wl[8302], wl[8303], wl[8304], wl[8305], wl[8306], wl[8307], wl[8308], wl[8309], wl[8310], wl[8311], wl[8312], wl[8313], wl[8314], wl[8315], wl[8316], wl[8317], wl[8318], wl[8319], wl[8320], wl[8321], wl[8322], wl[8323], wl[8324], wl[8325], wl[8326], wl[8327], wl[8328], wl[8329], wl[8330], wl[8331], wl[8332], wl[8333], wl[8334], wl[8335], wl[8336], wl[8337], wl[8338], wl[8339], wl[8340], wl[8341], wl[8342], wl[8343], wl[8344], wl[8345], wl[8346], wl[8347], wl[8348], wl[8349], wl[8350], wl[8351], wl[8352], wl[8353], wl[8354], wl[8355], wl[8356], wl[8357], wl[8358], wl[8359], wl[8360], wl[8361], wl[8362], wl[8363], wl[8364], wl[8365], wl[8366], wl[8367], wl[8368], wl[8369], wl[8370], wl[8371], wl[8372], wl[8373], wl[8374], wl[8375], wl[8376], wl[8377], wl[8378], wl[8379], wl[8380], wl[8381], wl[8382], wl[8383], wl[8384], wl[8385], wl[8386], wl[8387], wl[8388], wl[8389], wl[8390], wl[8391], wl[8392], wl[8393], wl[8394], wl[8395], wl[8396], wl[8397], wl[8398], wl[8399], wl[8400], wl[8401], wl[8402], wl[8403], wl[8404], wl[8405], wl[8406], wl[8407], wl[8408], wl[8409], wl[8410], wl[8411], wl[8412], wl[8413], wl[8414], wl[8415], wl[8416], wl[8417], wl[8418], wl[8419], wl[8420], wl[8421], wl[8422], wl[8423], wl[8424], wl[8425], wl[8426], wl[8427], wl[8428], wl[8429], wl[8430], wl[8431], wl[8432], wl[8433], wl[8434], wl[8435], wl[8436], wl[8437], wl[8438], wl[8439], wl[8440], wl[8441], wl[8442], wl[8443], wl[8444], wl[8445], wl[8446], wl[8447], wl[8448], wl[8449], wl[8450], wl[8451], wl[8452], wl[8453], wl[8454], wl[8455], wl[8456], wl[8457], wl[8458], wl[8459], wl[8460], wl[8461], wl[8462], wl[8463], wl[8464], wl[8465], wl[8466], wl[8467], wl[8468], wl[8469], wl[8470], wl[8471], wl[8472], wl[8473], wl[8474], wl[8475], wl[8476], wl[8477], wl[8478], wl[8479], wl[8480], wl[8481], wl[8482], wl[8483], wl[8484], wl[8485], wl[8486], wl[8487], wl[8488], wl[8489], wl[8490], wl[8491], wl[8492], wl[8493], wl[8494], wl[8495], wl[8496], wl[8497], wl[8498], wl[8499], wl[8500], wl[8501], wl[8502], wl[8503], wl[8504], wl[8505], wl[8506], wl[8507], wl[8508], wl[8509], wl[8510], wl[8511], wl[8512], wl[8513], wl[8514], wl[8515], wl[8516], wl[8517], wl[8518], wl[8519], wl[8520], wl[8521], wl[8522], wl[8523], wl[8524], wl[8525], wl[8526], wl[8527], wl[8528], wl[8529], wl[8530], wl[8531], wl[8532], wl[8533], wl[8534], wl[8535], wl[8536], wl[8537], wl[8538], wl[8539], wl[8540], wl[8541], wl[8542], wl[8543], wl[8544], wl[8545], wl[8546], wl[8547], wl[8548], wl[8549], wl[8550], wl[8551], wl[8552], wl[8553], wl[8554], wl[8555], wl[8556], wl[8557], wl[8558], wl[8559], wl[8560], wl[8561], wl[8562], wl[8563], wl[8564], wl[8565], wl[8566], wl[8567], wl[8568], wl[8569], wl[8570], wl[8571], wl[8572], wl[8573], wl[8574], wl[8575], wl[8576], wl[8577], wl[8578], wl[8579], wl[8580], wl[8581], wl[8582], wl[8583], wl[8584], wl[8585], wl[8586], wl[8587], wl[8588], wl[8589], wl[8590], wl[8591], wl[8592], wl[8593], wl[8594], wl[8595], wl[8596], wl[8597], wl[8598], wl[8599], wl[8600], wl[8601], wl[8602], wl[8603], wl[8604], wl[8605], wl[8606], wl[8607], wl[8608], wl[8609], wl[8610], wl[8611], wl[8612], wl[8613], wl[8614], wl[8615], wl[8616], wl[8617], wl[8618], wl[8619], wl[8620], wl[8621], wl[8622], wl[8623], wl[8624], wl[8625], wl[8626], wl[8627], wl[8628], wl[8629], wl[8630], wl[8631], wl[8632], wl[8633], wl[8634], wl[8635], wl[8636], wl[8637], wl[8638], wl[8639], wl[8640], wl[8641], wl[8642], wl[8643], wl[8644], wl[8645], wl[8646], wl[8647], wl[8648], wl[8649], wl[8650], wl[8651], wl[8652], wl[8653], wl[8654], wl[8655], wl[8656], wl[8657], wl[8658], wl[8659], wl[8660], wl[8661], wl[8662], wl[8663], wl[8664], wl[8665], wl[8666], wl[8667], wl[8668], wl[8669], wl[8670], wl[8671], wl[8672], wl[8673], wl[8674], wl[8675], wl[8676], wl[8677], wl[8678], wl[8679], wl[8680], wl[8681], wl[8682], wl[8683], wl[8684], wl[8685], wl[8686], wl[8687], wl[8688], wl[8689], wl[8690], wl[8691], wl[8692], wl[8693], wl[8694], wl[8695], wl[8696], wl[8697], wl[8698], wl[8699], wl[8700], wl[8701], wl[8702], wl[8703], wl[8704], wl[8705], wl[8706], wl[8707], wl[8708], wl[8709], wl[8710], wl[8711], wl[8712], wl[8713], wl[8714], wl[8715], wl[8716], wl[8717], wl[8718], wl[8719], wl[8720], wl[8721], wl[8722], wl[8723], wl[8724], wl[8725], wl[8726], wl[8727], wl[8728], wl[8729], wl[8730], wl[8731], wl[8732], wl[8733], wl[8734], wl[8735], wl[8736], wl[8737], wl[8738], wl[8739], wl[8740], wl[8741], wl[8742], wl[8743], wl[8744], wl[8745], wl[8746], wl[8747], wl[8748], wl[8749], wl[8750], wl[8751], wl[8752], wl[8753], wl[8754], wl[8755], wl[8756], wl[8757], wl[8758], wl[8759], wl[8760], wl[8761], wl[8762], wl[8763], wl[8764], wl[8765], wl[8766], wl[8767], wl[8768], wl[8769], wl[8770], wl[8771], wl[8772], wl[8773], wl[8774], wl[8775], wl[8776], wl[8777], wl[8778], wl[8779], wl[8780], wl[8781], wl[8782], wl[8783], wl[8784], wl[8785], wl[8786], wl[8787], wl[8788], wl[8789], wl[8790], wl[8791], wl[8792], wl[8793], wl[8794], wl[8795], wl[8796], wl[8797], wl[8798], wl[8799], wl[8800], wl[8801], wl[8802], wl[8803], wl[8804], wl[8805], wl[8806], wl[8807], wl[8808], wl[8809], wl[8810], wl[8811], wl[8812], wl[8813], wl[8814], wl[8815], wl[8816], wl[8817], wl[8818], wl[8819], wl[8820], wl[8821], wl[8822], wl[8823], wl[8824], wl[8825], wl[8826], wl[8827], wl[8828], wl[8829], wl[8830], wl[8831], wl[8832], wl[8833], wl[8834], wl[8835], wl[8836], wl[8837], wl[8838], wl[8839], wl[8840], wl[8841], wl[8842], wl[8843], wl[8844], wl[8845], wl[8846], wl[8847], wl[8848], wl[8849], wl[8850], wl[8851], wl[8852], wl[8853], wl[8854], wl[8855], wl[8856], wl[8857], wl[8858], wl[8859], wl[8860], wl[8861], wl[8862], wl[8863], wl[8864], wl[8865], wl[8866], wl[8867], wl[8868], wl[8869], wl[8870], wl[8871], wl[8872], wl[8873], wl[8874], wl[8875], wl[8876], wl[8877], wl[8878], wl[8879], wl[8880], wl[8881], wl[8882], wl[8883], wl[8884], wl[8885], wl[8886], wl[8887], wl[8888], wl[8889], wl[8890], wl[8891], wl[8892], wl[8893], wl[8894], wl[8895], wl[8896], wl[8897], wl[8898], wl[8899], wl[8900], wl[8901], wl[8902], wl[8903], wl[8904], wl[8905], wl[8906], wl[8907], wl[8908], wl[8909], wl[8910], wl[8911], wl[8912], wl[8913], wl[8914], wl[8915], wl[8916], wl[8917], wl[8918], wl[8919], wl[8920], wl[8921], wl[8922], wl[8923], wl[14044], wl[14045], wl[14046], wl[14047], wl[14048], wl[14049], wl[14050], wl[14051], wl[14052], wl[14053], wl[14054], wl[14055], wl[14056], wl[14057], wl[14058], wl[14059], wl[14060], wl[14061], wl[14062], wl[14063], wl[14064], wl[14065], wl[14066], wl[14067], wl[14068], wl[14069], wl[14070], wl[14071], wl[14072], wl[14073], wl[14074], wl[14075], wl[14076], wl[14077], wl[14078], wl[14079], wl[14080], wl[14081], wl[14082], wl[14083], wl[14084], wl[14085], wl[14086], wl[14087], wl[14088], wl[14089], wl[14090], wl[14091], wl[14092], wl[14093], wl[14094], wl[14095], wl[14096], wl[14097], wl[14098], wl[14099], wl[14100], wl[14101], wl[14102], wl[14103], wl[14104], wl[14105], wl[14106], wl[14107], wl[14108], wl[14109], wl[14110], wl[14111], wl[14112], wl[14113], wl[14114], wl[14115], wl[14116], wl[14117], wl[14118], wl[14119], wl[14120], wl[14121], wl[14122], wl[14123], wl[7824], wl[7825], wl[7826], wl[7827], wl[7828], wl[7829], wl[7830], wl[7831], wl[7832], wl[7833], wl[7834], wl[7835], wl[7836], wl[7837], wl[7838], wl[7839], wl[7840], wl[7841], wl[7842], wl[7843], wl[7844], wl[7845], wl[7846], wl[7847], wl[7848], wl[7849], wl[7850], wl[7851], wl[7852], wl[7853], wl[7854], wl[7855], wl[7856], wl[7857], wl[7858], wl[7859], wl[7860], wl[7861], wl[7862], wl[7863], wl[7864], wl[7865], wl[7866], wl[7867], wl[7868], wl[7869], wl[7870], wl[7871], wl[7872], wl[7873], wl[7874], wl[7875], wl[7876], wl[7877], wl[7878], wl[7879], wl[7880], wl[7881], wl[7882], wl[7883], wl[7884], wl[7885], wl[7886], wl[7887], wl[7888], wl[7889], wl[7890], wl[7891], wl[7892], wl[7893], wl[7894], wl[7895], wl[7896], wl[7897], wl[7898], wl[7899], wl[7900], wl[7901], wl[7902], wl[7903], wl[13964], wl[13965], wl[13966], wl[13967], wl[13968], wl[13969], wl[13970], wl[13971], wl[13972], wl[13973], wl[13974], wl[13975], wl[13976], wl[13977], wl[13978], wl[13979], wl[13980], wl[13981], wl[13982], wl[13983], wl[13984], wl[13985], wl[13986], wl[13987], wl[13988], wl[13989], wl[13990], wl[13991], wl[13992], wl[13993], wl[13994], wl[13995], wl[13996], wl[13997], wl[13998], wl[13999], wl[14000], wl[14001], wl[14002], wl[14003], wl[14004], wl[14005], wl[14006], wl[14007], wl[14008], wl[14009], wl[14010], wl[14011], wl[14012], wl[14013], wl[14014], wl[14015], wl[14016], wl[14017], wl[14018], wl[14019], wl[14020], wl[14021], wl[14022], wl[14023], wl[14024], wl[14025], wl[14026], wl[14027], wl[14028], wl[14029], wl[14030], wl[14031], wl[14032], wl[14033], wl[14034], wl[14035], wl[14036], wl[14037], wl[14038], wl[14039], wl[14040], wl[14041], wl[14042], wl[14043]})
    );
    tile tile_4__4_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_2__3__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_2__3__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_2__3__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_3__2__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_3__2__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_3__2__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_2__2__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_2__2__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_2__2__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_2__2__grid_top_r_in[1]),
        .grid_left_in(grid_clb_3__3__grid_left_in),
        .grid_bottom_in(grid_clb_3__3__grid_bottom_in),
        .chanx_left_in(sb_1__1__5_chanx_right_out),
        .chanx_left_out(cbx_1__1__8_chanx_left_out),
        .grid_top_out(grid_clb_3__4__grid_bottom_in),
        .chany_bottom_in(sb_1__1__7_chany_top_out),
        .chany_bottom_out(cby_1__1__10_chany_bottom_out),
        .grid_right_out(grid_clb_4__3__grid_left_in),
        .chany_top_in_0(cby_1__1__11_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__11_chanx_left_out),
        .chany_top_out_0(sb_1__1__8_chany_top_out),
        .chanx_right_out_0(sb_1__1__8_chanx_right_out),
        .grid_top_r_in(sb_3__3__grid_top_r_in),
        .grid_top_l_in(sb_3__3__grid_top_l_in),
        .grid_right_t_in(sb_3__3__grid_right_t_in),
        .grid_right_b_in(sb_3__3__grid_right_b_in),
        .grid_bottom_r_in(sb_3__2__grid_top_r_in),
        .grid_bottom_l_in(sb_3__2__grid_top_l_in),
        .grid_left_t_in(sb_2__3__grid_right_t_in),
        .grid_left_b_in(sb_2__3__grid_right_b_in),
        .bl({bl[14204], bl[14205], bl[14206], bl[14207], bl[14208], bl[14209], bl[14210], bl[14211], bl[14212], bl[14213], bl[14214], bl[14215], bl[14216], bl[14217], bl[14218], bl[14219], bl[14220], bl[14221], bl[14222], bl[14223], bl[14224], bl[14225], bl[14226], bl[14227], bl[14228], bl[14229], bl[14230], bl[14231], bl[14232], bl[14233], bl[14234], bl[14235], bl[14236], bl[14237], bl[14238], bl[14239], bl[14240], bl[14241], bl[14242], bl[14243], bl[14244], bl[14245], bl[14246], bl[14247], bl[14248], bl[14249], bl[14250], bl[14251], bl[14252], bl[14253], bl[14254], bl[14255], bl[14256], bl[14257], bl[14258], bl[14259], bl[14260], bl[14261], bl[14262], bl[14263], bl[14264], bl[14265], bl[14266], bl[14267], bl[14268], bl[14269], bl[14270], bl[14271], bl[14272], bl[14273], bl[14274], bl[14275], bl[14276], bl[14277], bl[14278], bl[14279], bl[14280], bl[14281], bl[14282], bl[14283], bl[14284], bl[14285], bl[14286], bl[14287], bl[14288], bl[14289], bl[14290], bl[14291], bl[14292], bl[14293], bl[14294], bl[14295], bl[14296], bl[14297], bl[14298], bl[14299], bl[14300], bl[14301], bl[14302], bl[14303], bl[14304], bl[14305], bl[14306], bl[14307], bl[14308], bl[14309], bl[14310], bl[14311], bl[14312], bl[14313], bl[14314], bl[14315], bl[14316], bl[14317], bl[14318], bl[14319], bl[14320], bl[14321], bl[14322], bl[14323], bl[14324], bl[14325], bl[14326], bl[14327], bl[14328], bl[14329], bl[14330], bl[14331], bl[14332], bl[14333], bl[14334], bl[14335], bl[14336], bl[14337], bl[14338], bl[14339], bl[14340], bl[14341], bl[14342], bl[14343], bl[14344], bl[14345], bl[14346], bl[14347], bl[14348], bl[14349], bl[14350], bl[14351], bl[14352], bl[14353], bl[14354], bl[14355], bl[14356], bl[14357], bl[14358], bl[14359], bl[14360], bl[14361], bl[14362], bl[14363], bl[14364], bl[14365], bl[14366], bl[14367], bl[14368], bl[14369], bl[14370], bl[14371], bl[14372], bl[14373], bl[14374], bl[14375], bl[14376], bl[14377], bl[14378], bl[14379], bl[14380], bl[14381], bl[14382], bl[14383], bl[14384], bl[14385], bl[14386], bl[14387], bl[14388], bl[14389], bl[14390], bl[14391], bl[14392], bl[14393], bl[14394], bl[14395], bl[14396], bl[14397], bl[14398], bl[14399], bl[14400], bl[14401], bl[14402], bl[14403], bl[14404], bl[14405], bl[14406], bl[14407], bl[14408], bl[14409], bl[14410], bl[14411], bl[14412], bl[14413], bl[14414], bl[14415], bl[14416], bl[14417], bl[14418], bl[14419], bl[14420], bl[14421], bl[14422], bl[14423], bl[14424], bl[14425], bl[14426], bl[14427], bl[14428], bl[14429], bl[14430], bl[14431], bl[14432], bl[14433], bl[14434], bl[14435], bl[14436], bl[14437], bl[14438], bl[14439], bl[14440], bl[14441], bl[14442], bl[14443], bl[14444], bl[14445], bl[14446], bl[14447], bl[14448], bl[14449], bl[14450], bl[14451], bl[14452], bl[14453], bl[14454], bl[14455], bl[14456], bl[14457], bl[14458], bl[14459], bl[14460], bl[14461], bl[14462], bl[14463], bl[14464], bl[14465], bl[14466], bl[14467], bl[14468], bl[14469], bl[14470], bl[14471], bl[14472], bl[14473], bl[14474], bl[14475], bl[14476], bl[14477], bl[14478], bl[14479], bl[14480], bl[14481], bl[14482], bl[14483], bl[14484], bl[14485], bl[14486], bl[14487], bl[14488], bl[14489], bl[14490], bl[14491], bl[14492], bl[14493], bl[14494], bl[14495], bl[14496], bl[14497], bl[14498], bl[14499], bl[14500], bl[14501], bl[14502], bl[14503], bl[14504], bl[14505], bl[14506], bl[14507], bl[14508], bl[14509], bl[14510], bl[14511], bl[14512], bl[14513], bl[14514], bl[14515], bl[14516], bl[14517], bl[14518], bl[14519], bl[14520], bl[14521], bl[14522], bl[14523], bl[14524], bl[14525], bl[14526], bl[14527], bl[14528], bl[14529], bl[14530], bl[14531], bl[14532], bl[14533], bl[14534], bl[14535], bl[14536], bl[14537], bl[14538], bl[14539], bl[14540], bl[14541], bl[14542], bl[14543], bl[14544], bl[14545], bl[14546], bl[14547], bl[14548], bl[14549], bl[14550], bl[14551], bl[14552], bl[14553], bl[14554], bl[14555], bl[14556], bl[14557], bl[14558], bl[14559], bl[14560], bl[14561], bl[14562], bl[14563], bl[14564], bl[14565], bl[14566], bl[14567], bl[14568], bl[14569], bl[14570], bl[14571], bl[14572], bl[14573], bl[14574], bl[14575], bl[14576], bl[14577], bl[14578], bl[14579], bl[14580], bl[14581], bl[14582], bl[14583], bl[14584], bl[14585], bl[14586], bl[14587], bl[14588], bl[14589], bl[14590], bl[14591], bl[14592], bl[14593], bl[14594], bl[14595], bl[14596], bl[14597], bl[14598], bl[14599], bl[14600], bl[14601], bl[14602], bl[14603], bl[14604], bl[14605], bl[14606], bl[14607], bl[14608], bl[14609], bl[14610], bl[14611], bl[14612], bl[14613], bl[14614], bl[14615], bl[14616], bl[14617], bl[14618], bl[14619], bl[14620], bl[14621], bl[14622], bl[14623], bl[14624], bl[14625], bl[14626], bl[14627], bl[14628], bl[14629], bl[14630], bl[14631], bl[14632], bl[14633], bl[14634], bl[14635], bl[14636], bl[14637], bl[14638], bl[14639], bl[14640], bl[14641], bl[14642], bl[14643], bl[14644], bl[14645], bl[14646], bl[14647], bl[14648], bl[14649], bl[14650], bl[14651], bl[14652], bl[14653], bl[14654], bl[14655], bl[14656], bl[14657], bl[14658], bl[14659], bl[14660], bl[14661], bl[14662], bl[14663], bl[14664], bl[14665], bl[14666], bl[14667], bl[14668], bl[14669], bl[14670], bl[14671], bl[14672], bl[14673], bl[14674], bl[14675], bl[14676], bl[14677], bl[14678], bl[14679], bl[14680], bl[14681], bl[14682], bl[14683], bl[14684], bl[14685], bl[14686], bl[14687], bl[14688], bl[14689], bl[14690], bl[14691], bl[14692], bl[14693], bl[14694], bl[14695], bl[14696], bl[14697], bl[14698], bl[14699], bl[14700], bl[14701], bl[14702], bl[14703], bl[14704], bl[14705], bl[14706], bl[14707], bl[14708], bl[14709], bl[14710], bl[14711], bl[14712], bl[14713], bl[14714], bl[14715], bl[14716], bl[14717], bl[14718], bl[14719], bl[14720], bl[14721], bl[14722], bl[14723], bl[14724], bl[14725], bl[14726], bl[14727], bl[14728], bl[14729], bl[14730], bl[14731], bl[14732], bl[14733], bl[14734], bl[14735], bl[14736], bl[14737], bl[14738], bl[14739], bl[14740], bl[14741], bl[14742], bl[14743], bl[14744], bl[14745], bl[14746], bl[14747], bl[14748], bl[14749], bl[14750], bl[14751], bl[14752], bl[14753], bl[14754], bl[14755], bl[14756], bl[14757], bl[14758], bl[14759], bl[14760], bl[14761], bl[14762], bl[14763], bl[14764], bl[14765], bl[14766], bl[14767], bl[14768], bl[14769], bl[14770], bl[14771], bl[14772], bl[14773], bl[14774], bl[14775], bl[14776], bl[14777], bl[14778], bl[14779], bl[14780], bl[14781], bl[14782], bl[14783], bl[14784], bl[14785], bl[14786], bl[14787], bl[14788], bl[14789], bl[14790], bl[14791], bl[14792], bl[14793], bl[14794], bl[14795], bl[14796], bl[14797], bl[14798], bl[14799], bl[14800], bl[14801], bl[14802], bl[14803], bl[14804], bl[14805], bl[14806], bl[14807], bl[14808], bl[14809], bl[14810], bl[14811], bl[14812], bl[14813], bl[14814], bl[14815], bl[14816], bl[14817], bl[14818], bl[14819], bl[14820], bl[14821], bl[14822], bl[14823], bl[14824], bl[14825], bl[14826], bl[14827], bl[14828], bl[14829], bl[14830], bl[14831], bl[14832], bl[14833], bl[14834], bl[14835], bl[14836], bl[14837], bl[14838], bl[14839], bl[14840], bl[14841], bl[14842], bl[14843], bl[14844], bl[14845], bl[14846], bl[14847], bl[14848], bl[14849], bl[14850], bl[14851], bl[14852], bl[14853], bl[14854], bl[14855], bl[14856], bl[14857], bl[14858], bl[14859], bl[14860], bl[14861], bl[14862], bl[14863], bl[14864], bl[14865], bl[14866], bl[14867], bl[14868], bl[14869], bl[14870], bl[14871], bl[14872], bl[14873], bl[14874], bl[14875], bl[14876], bl[14877], bl[14878], bl[14879], bl[14880], bl[14881], bl[14882], bl[14883], bl[14884], bl[14885], bl[14886], bl[14887], bl[14888], bl[14889], bl[14890], bl[14891], bl[14892], bl[14893], bl[14894], bl[14895], bl[14896], bl[14897], bl[14898], bl[14899], bl[14900], bl[14901], bl[14902], bl[14903], bl[14904], bl[14905], bl[14906], bl[14907], bl[14908], bl[14909], bl[14910], bl[14911], bl[14912], bl[14913], bl[14914], bl[14915], bl[14916], bl[14917], bl[14918], bl[14919], bl[14920], bl[14921], bl[14922], bl[14923], bl[14924], bl[14925], bl[14926], bl[14927], bl[14928], bl[14929], bl[14930], bl[14931], bl[14932], bl[14933], bl[14934], bl[14935], bl[14936], bl[14937], bl[14938], bl[14939], bl[14940], bl[14941], bl[14942], bl[14943], bl[14944], bl[14945], bl[14946], bl[14947], bl[14948], bl[14949], bl[14950], bl[14951], bl[14952], bl[14953], bl[14954], bl[14955], bl[14956], bl[14957], bl[14958], bl[14959], bl[14960], bl[14961], bl[14962], bl[14963], bl[14964], bl[14965], bl[14966], bl[14967], bl[14968], bl[14969], bl[14970], bl[14971], bl[14972], bl[14973], bl[14974], bl[14975], bl[14976], bl[14977], bl[14978], bl[14979], bl[14980], bl[14981], bl[14982], bl[14983], bl[14984], bl[14985], bl[14986], bl[14987], bl[14988], bl[14989], bl[14990], bl[14991], bl[14992], bl[14993], bl[14994], bl[14995], bl[14996], bl[14997], bl[14998], bl[14999], bl[15000], bl[15001], bl[15002], bl[15003], bl[15004], bl[15005], bl[15006], bl[15007], bl[15008], bl[15009], bl[15010], bl[15011], bl[15012], bl[15013], bl[15014], bl[15015], bl[15016], bl[15017], bl[15018], bl[15019], bl[15020], bl[15021], bl[15022], bl[15023], bl[15024], bl[15025], bl[15026], bl[15027], bl[15028], bl[15029], bl[15030], bl[15031], bl[15032], bl[15033], bl[15034], bl[15035], bl[15036], bl[15037], bl[15038], bl[15039], bl[15040], bl[15041], bl[15042], bl[15043], bl[15044], bl[15045], bl[15046], bl[15047], bl[15048], bl[15049], bl[15050], bl[15051], bl[15052], bl[15053], bl[15054], bl[15055], bl[15056], bl[15057], bl[15058], bl[15059], bl[15060], bl[15061], bl[15062], bl[15063], bl[15064], bl[15065], bl[15066], bl[15067], bl[15068], bl[15069], bl[15070], bl[15071], bl[15072], bl[15073], bl[15074], bl[15075], bl[15076], bl[15077], bl[15078], bl[15079], bl[15080], bl[15081], bl[15082], bl[15083], bl[15084], bl[15085], bl[15086], bl[15087], bl[15088], bl[15089], bl[15090], bl[15091], bl[15092], bl[15093], bl[15094], bl[15095], bl[15096], bl[15097], bl[15098], bl[15099], bl[15100], bl[15101], bl[15102], bl[15103], bl[15104], bl[15105], bl[15106], bl[15107], bl[15108], bl[15109], bl[15110], bl[15111], bl[15112], bl[15113], bl[15114], bl[15115], bl[15116], bl[15117], bl[15118], bl[15119], bl[15120], bl[15121], bl[15122], bl[15123], bl[15124], bl[15125], bl[15126], bl[15127], bl[15128], bl[15129], bl[15130], bl[15131], bl[15132], bl[15133], bl[15134], bl[15135], bl[15136], bl[15137], bl[15138], bl[15139], bl[15140], bl[15141], bl[15142], bl[15143], bl[15144], bl[15145], bl[15146], bl[15147], bl[15148], bl[15149], bl[15150], bl[15151], bl[15152], bl[15153], bl[15154], bl[15155], bl[15156], bl[15157], bl[15158], bl[15159], bl[15160], bl[15161], bl[15162], bl[15163], bl[15164], bl[15165], bl[15166], bl[15167], bl[15168], bl[15169], bl[15170], bl[15171], bl[15172], bl[15173], bl[15174], bl[15175], bl[15176], bl[15177], bl[15178], bl[15179], bl[15180], bl[15181], bl[15182], bl[15183], bl[15184], bl[15185], bl[15186], bl[15187], bl[15188], bl[15189], bl[15190], bl[15191], bl[15192], bl[15193], bl[15194], bl[15195], bl[15196], bl[15197], bl[15198], bl[15199], bl[15200], bl[15201], bl[15202], bl[15203], bl[15204], bl[15205], bl[15206], bl[15207], bl[15208], bl[15209], bl[15210], bl[15211], bl[15212], bl[15213], bl[15214], bl[15215], bl[15216], bl[15217], bl[15218], bl[15219], bl[15220], bl[15221], bl[15222], bl[15223], bl[17808], bl[17809], bl[17810], bl[17811], bl[17812], bl[17813], bl[17814], bl[17815], bl[17816], bl[17817], bl[17818], bl[17819], bl[17820], bl[17821], bl[17822], bl[17823], bl[17824], bl[17825], bl[17826], bl[17827], bl[17828], bl[17829], bl[17830], bl[17831], bl[17832], bl[17833], bl[17834], bl[17835], bl[17836], bl[17837], bl[17838], bl[17839], bl[17840], bl[17841], bl[17842], bl[17843], bl[17844], bl[17845], bl[17846], bl[17847], bl[17848], bl[17849], bl[17850], bl[17851], bl[17852], bl[17853], bl[17854], bl[17855], bl[17856], bl[17857], bl[17858], bl[17859], bl[17860], bl[17861], bl[17862], bl[17863], bl[17864], bl[17865], bl[17866], bl[17867], bl[17868], bl[17869], bl[17870], bl[17871], bl[17872], bl[17873], bl[17874], bl[17875], bl[17876], bl[17877], bl[17878], bl[17879], bl[17880], bl[17881], bl[17882], bl[17883], bl[17884], bl[17885], bl[17886], bl[17887], bl[14124], bl[14125], bl[14126], bl[14127], bl[14128], bl[14129], bl[14130], bl[14131], bl[14132], bl[14133], bl[14134], bl[14135], bl[14136], bl[14137], bl[14138], bl[14139], bl[14140], bl[14141], bl[14142], bl[14143], bl[14144], bl[14145], bl[14146], bl[14147], bl[14148], bl[14149], bl[14150], bl[14151], bl[14152], bl[14153], bl[14154], bl[14155], bl[14156], bl[14157], bl[14158], bl[14159], bl[14160], bl[14161], bl[14162], bl[14163], bl[14164], bl[14165], bl[14166], bl[14167], bl[14168], bl[14169], bl[14170], bl[14171], bl[14172], bl[14173], bl[14174], bl[14175], bl[14176], bl[14177], bl[14178], bl[14179], bl[14180], bl[14181], bl[14182], bl[14183], bl[14184], bl[14185], bl[14186], bl[14187], bl[14188], bl[14189], bl[14190], bl[14191], bl[14192], bl[14193], bl[14194], bl[14195], bl[14196], bl[14197], bl[14198], bl[14199], bl[14200], bl[14201], bl[14202], bl[14203], bl[17728], bl[17729], bl[17730], bl[17731], bl[17732], bl[17733], bl[17734], bl[17735], bl[17736], bl[17737], bl[17738], bl[17739], bl[17740], bl[17741], bl[17742], bl[17743], bl[17744], bl[17745], bl[17746], bl[17747], bl[17748], bl[17749], bl[17750], bl[17751], bl[17752], bl[17753], bl[17754], bl[17755], bl[17756], bl[17757], bl[17758], bl[17759], bl[17760], bl[17761], bl[17762], bl[17763], bl[17764], bl[17765], bl[17766], bl[17767], bl[17768], bl[17769], bl[17770], bl[17771], bl[17772], bl[17773], bl[17774], bl[17775], bl[17776], bl[17777], bl[17778], bl[17779], bl[17780], bl[17781], bl[17782], bl[17783], bl[17784], bl[17785], bl[17786], bl[17787], bl[17788], bl[17789], bl[17790], bl[17791], bl[17792], bl[17793], bl[17794], bl[17795], bl[17796], bl[17797], bl[17798], bl[17799], bl[17800], bl[17801], bl[17802], bl[17803], bl[17804], bl[17805], bl[17806], bl[17807]}),
        .wl({wl[14204], wl[14205], wl[14206], wl[14207], wl[14208], wl[14209], wl[14210], wl[14211], wl[14212], wl[14213], wl[14214], wl[14215], wl[14216], wl[14217], wl[14218], wl[14219], wl[14220], wl[14221], wl[14222], wl[14223], wl[14224], wl[14225], wl[14226], wl[14227], wl[14228], wl[14229], wl[14230], wl[14231], wl[14232], wl[14233], wl[14234], wl[14235], wl[14236], wl[14237], wl[14238], wl[14239], wl[14240], wl[14241], wl[14242], wl[14243], wl[14244], wl[14245], wl[14246], wl[14247], wl[14248], wl[14249], wl[14250], wl[14251], wl[14252], wl[14253], wl[14254], wl[14255], wl[14256], wl[14257], wl[14258], wl[14259], wl[14260], wl[14261], wl[14262], wl[14263], wl[14264], wl[14265], wl[14266], wl[14267], wl[14268], wl[14269], wl[14270], wl[14271], wl[14272], wl[14273], wl[14274], wl[14275], wl[14276], wl[14277], wl[14278], wl[14279], wl[14280], wl[14281], wl[14282], wl[14283], wl[14284], wl[14285], wl[14286], wl[14287], wl[14288], wl[14289], wl[14290], wl[14291], wl[14292], wl[14293], wl[14294], wl[14295], wl[14296], wl[14297], wl[14298], wl[14299], wl[14300], wl[14301], wl[14302], wl[14303], wl[14304], wl[14305], wl[14306], wl[14307], wl[14308], wl[14309], wl[14310], wl[14311], wl[14312], wl[14313], wl[14314], wl[14315], wl[14316], wl[14317], wl[14318], wl[14319], wl[14320], wl[14321], wl[14322], wl[14323], wl[14324], wl[14325], wl[14326], wl[14327], wl[14328], wl[14329], wl[14330], wl[14331], wl[14332], wl[14333], wl[14334], wl[14335], wl[14336], wl[14337], wl[14338], wl[14339], wl[14340], wl[14341], wl[14342], wl[14343], wl[14344], wl[14345], wl[14346], wl[14347], wl[14348], wl[14349], wl[14350], wl[14351], wl[14352], wl[14353], wl[14354], wl[14355], wl[14356], wl[14357], wl[14358], wl[14359], wl[14360], wl[14361], wl[14362], wl[14363], wl[14364], wl[14365], wl[14366], wl[14367], wl[14368], wl[14369], wl[14370], wl[14371], wl[14372], wl[14373], wl[14374], wl[14375], wl[14376], wl[14377], wl[14378], wl[14379], wl[14380], wl[14381], wl[14382], wl[14383], wl[14384], wl[14385], wl[14386], wl[14387], wl[14388], wl[14389], wl[14390], wl[14391], wl[14392], wl[14393], wl[14394], wl[14395], wl[14396], wl[14397], wl[14398], wl[14399], wl[14400], wl[14401], wl[14402], wl[14403], wl[14404], wl[14405], wl[14406], wl[14407], wl[14408], wl[14409], wl[14410], wl[14411], wl[14412], wl[14413], wl[14414], wl[14415], wl[14416], wl[14417], wl[14418], wl[14419], wl[14420], wl[14421], wl[14422], wl[14423], wl[14424], wl[14425], wl[14426], wl[14427], wl[14428], wl[14429], wl[14430], wl[14431], wl[14432], wl[14433], wl[14434], wl[14435], wl[14436], wl[14437], wl[14438], wl[14439], wl[14440], wl[14441], wl[14442], wl[14443], wl[14444], wl[14445], wl[14446], wl[14447], wl[14448], wl[14449], wl[14450], wl[14451], wl[14452], wl[14453], wl[14454], wl[14455], wl[14456], wl[14457], wl[14458], wl[14459], wl[14460], wl[14461], wl[14462], wl[14463], wl[14464], wl[14465], wl[14466], wl[14467], wl[14468], wl[14469], wl[14470], wl[14471], wl[14472], wl[14473], wl[14474], wl[14475], wl[14476], wl[14477], wl[14478], wl[14479], wl[14480], wl[14481], wl[14482], wl[14483], wl[14484], wl[14485], wl[14486], wl[14487], wl[14488], wl[14489], wl[14490], wl[14491], wl[14492], wl[14493], wl[14494], wl[14495], wl[14496], wl[14497], wl[14498], wl[14499], wl[14500], wl[14501], wl[14502], wl[14503], wl[14504], wl[14505], wl[14506], wl[14507], wl[14508], wl[14509], wl[14510], wl[14511], wl[14512], wl[14513], wl[14514], wl[14515], wl[14516], wl[14517], wl[14518], wl[14519], wl[14520], wl[14521], wl[14522], wl[14523], wl[14524], wl[14525], wl[14526], wl[14527], wl[14528], wl[14529], wl[14530], wl[14531], wl[14532], wl[14533], wl[14534], wl[14535], wl[14536], wl[14537], wl[14538], wl[14539], wl[14540], wl[14541], wl[14542], wl[14543], wl[14544], wl[14545], wl[14546], wl[14547], wl[14548], wl[14549], wl[14550], wl[14551], wl[14552], wl[14553], wl[14554], wl[14555], wl[14556], wl[14557], wl[14558], wl[14559], wl[14560], wl[14561], wl[14562], wl[14563], wl[14564], wl[14565], wl[14566], wl[14567], wl[14568], wl[14569], wl[14570], wl[14571], wl[14572], wl[14573], wl[14574], wl[14575], wl[14576], wl[14577], wl[14578], wl[14579], wl[14580], wl[14581], wl[14582], wl[14583], wl[14584], wl[14585], wl[14586], wl[14587], wl[14588], wl[14589], wl[14590], wl[14591], wl[14592], wl[14593], wl[14594], wl[14595], wl[14596], wl[14597], wl[14598], wl[14599], wl[14600], wl[14601], wl[14602], wl[14603], wl[14604], wl[14605], wl[14606], wl[14607], wl[14608], wl[14609], wl[14610], wl[14611], wl[14612], wl[14613], wl[14614], wl[14615], wl[14616], wl[14617], wl[14618], wl[14619], wl[14620], wl[14621], wl[14622], wl[14623], wl[14624], wl[14625], wl[14626], wl[14627], wl[14628], wl[14629], wl[14630], wl[14631], wl[14632], wl[14633], wl[14634], wl[14635], wl[14636], wl[14637], wl[14638], wl[14639], wl[14640], wl[14641], wl[14642], wl[14643], wl[14644], wl[14645], wl[14646], wl[14647], wl[14648], wl[14649], wl[14650], wl[14651], wl[14652], wl[14653], wl[14654], wl[14655], wl[14656], wl[14657], wl[14658], wl[14659], wl[14660], wl[14661], wl[14662], wl[14663], wl[14664], wl[14665], wl[14666], wl[14667], wl[14668], wl[14669], wl[14670], wl[14671], wl[14672], wl[14673], wl[14674], wl[14675], wl[14676], wl[14677], wl[14678], wl[14679], wl[14680], wl[14681], wl[14682], wl[14683], wl[14684], wl[14685], wl[14686], wl[14687], wl[14688], wl[14689], wl[14690], wl[14691], wl[14692], wl[14693], wl[14694], wl[14695], wl[14696], wl[14697], wl[14698], wl[14699], wl[14700], wl[14701], wl[14702], wl[14703], wl[14704], wl[14705], wl[14706], wl[14707], wl[14708], wl[14709], wl[14710], wl[14711], wl[14712], wl[14713], wl[14714], wl[14715], wl[14716], wl[14717], wl[14718], wl[14719], wl[14720], wl[14721], wl[14722], wl[14723], wl[14724], wl[14725], wl[14726], wl[14727], wl[14728], wl[14729], wl[14730], wl[14731], wl[14732], wl[14733], wl[14734], wl[14735], wl[14736], wl[14737], wl[14738], wl[14739], wl[14740], wl[14741], wl[14742], wl[14743], wl[14744], wl[14745], wl[14746], wl[14747], wl[14748], wl[14749], wl[14750], wl[14751], wl[14752], wl[14753], wl[14754], wl[14755], wl[14756], wl[14757], wl[14758], wl[14759], wl[14760], wl[14761], wl[14762], wl[14763], wl[14764], wl[14765], wl[14766], wl[14767], wl[14768], wl[14769], wl[14770], wl[14771], wl[14772], wl[14773], wl[14774], wl[14775], wl[14776], wl[14777], wl[14778], wl[14779], wl[14780], wl[14781], wl[14782], wl[14783], wl[14784], wl[14785], wl[14786], wl[14787], wl[14788], wl[14789], wl[14790], wl[14791], wl[14792], wl[14793], wl[14794], wl[14795], wl[14796], wl[14797], wl[14798], wl[14799], wl[14800], wl[14801], wl[14802], wl[14803], wl[14804], wl[14805], wl[14806], wl[14807], wl[14808], wl[14809], wl[14810], wl[14811], wl[14812], wl[14813], wl[14814], wl[14815], wl[14816], wl[14817], wl[14818], wl[14819], wl[14820], wl[14821], wl[14822], wl[14823], wl[14824], wl[14825], wl[14826], wl[14827], wl[14828], wl[14829], wl[14830], wl[14831], wl[14832], wl[14833], wl[14834], wl[14835], wl[14836], wl[14837], wl[14838], wl[14839], wl[14840], wl[14841], wl[14842], wl[14843], wl[14844], wl[14845], wl[14846], wl[14847], wl[14848], wl[14849], wl[14850], wl[14851], wl[14852], wl[14853], wl[14854], wl[14855], wl[14856], wl[14857], wl[14858], wl[14859], wl[14860], wl[14861], wl[14862], wl[14863], wl[14864], wl[14865], wl[14866], wl[14867], wl[14868], wl[14869], wl[14870], wl[14871], wl[14872], wl[14873], wl[14874], wl[14875], wl[14876], wl[14877], wl[14878], wl[14879], wl[14880], wl[14881], wl[14882], wl[14883], wl[14884], wl[14885], wl[14886], wl[14887], wl[14888], wl[14889], wl[14890], wl[14891], wl[14892], wl[14893], wl[14894], wl[14895], wl[14896], wl[14897], wl[14898], wl[14899], wl[14900], wl[14901], wl[14902], wl[14903], wl[14904], wl[14905], wl[14906], wl[14907], wl[14908], wl[14909], wl[14910], wl[14911], wl[14912], wl[14913], wl[14914], wl[14915], wl[14916], wl[14917], wl[14918], wl[14919], wl[14920], wl[14921], wl[14922], wl[14923], wl[14924], wl[14925], wl[14926], wl[14927], wl[14928], wl[14929], wl[14930], wl[14931], wl[14932], wl[14933], wl[14934], wl[14935], wl[14936], wl[14937], wl[14938], wl[14939], wl[14940], wl[14941], wl[14942], wl[14943], wl[14944], wl[14945], wl[14946], wl[14947], wl[14948], wl[14949], wl[14950], wl[14951], wl[14952], wl[14953], wl[14954], wl[14955], wl[14956], wl[14957], wl[14958], wl[14959], wl[14960], wl[14961], wl[14962], wl[14963], wl[14964], wl[14965], wl[14966], wl[14967], wl[14968], wl[14969], wl[14970], wl[14971], wl[14972], wl[14973], wl[14974], wl[14975], wl[14976], wl[14977], wl[14978], wl[14979], wl[14980], wl[14981], wl[14982], wl[14983], wl[14984], wl[14985], wl[14986], wl[14987], wl[14988], wl[14989], wl[14990], wl[14991], wl[14992], wl[14993], wl[14994], wl[14995], wl[14996], wl[14997], wl[14998], wl[14999], wl[15000], wl[15001], wl[15002], wl[15003], wl[15004], wl[15005], wl[15006], wl[15007], wl[15008], wl[15009], wl[15010], wl[15011], wl[15012], wl[15013], wl[15014], wl[15015], wl[15016], wl[15017], wl[15018], wl[15019], wl[15020], wl[15021], wl[15022], wl[15023], wl[15024], wl[15025], wl[15026], wl[15027], wl[15028], wl[15029], wl[15030], wl[15031], wl[15032], wl[15033], wl[15034], wl[15035], wl[15036], wl[15037], wl[15038], wl[15039], wl[15040], wl[15041], wl[15042], wl[15043], wl[15044], wl[15045], wl[15046], wl[15047], wl[15048], wl[15049], wl[15050], wl[15051], wl[15052], wl[15053], wl[15054], wl[15055], wl[15056], wl[15057], wl[15058], wl[15059], wl[15060], wl[15061], wl[15062], wl[15063], wl[15064], wl[15065], wl[15066], wl[15067], wl[15068], wl[15069], wl[15070], wl[15071], wl[15072], wl[15073], wl[15074], wl[15075], wl[15076], wl[15077], wl[15078], wl[15079], wl[15080], wl[15081], wl[15082], wl[15083], wl[15084], wl[15085], wl[15086], wl[15087], wl[15088], wl[15089], wl[15090], wl[15091], wl[15092], wl[15093], wl[15094], wl[15095], wl[15096], wl[15097], wl[15098], wl[15099], wl[15100], wl[15101], wl[15102], wl[15103], wl[15104], wl[15105], wl[15106], wl[15107], wl[15108], wl[15109], wl[15110], wl[15111], wl[15112], wl[15113], wl[15114], wl[15115], wl[15116], wl[15117], wl[15118], wl[15119], wl[15120], wl[15121], wl[15122], wl[15123], wl[15124], wl[15125], wl[15126], wl[15127], wl[15128], wl[15129], wl[15130], wl[15131], wl[15132], wl[15133], wl[15134], wl[15135], wl[15136], wl[15137], wl[15138], wl[15139], wl[15140], wl[15141], wl[15142], wl[15143], wl[15144], wl[15145], wl[15146], wl[15147], wl[15148], wl[15149], wl[15150], wl[15151], wl[15152], wl[15153], wl[15154], wl[15155], wl[15156], wl[15157], wl[15158], wl[15159], wl[15160], wl[15161], wl[15162], wl[15163], wl[15164], wl[15165], wl[15166], wl[15167], wl[15168], wl[15169], wl[15170], wl[15171], wl[15172], wl[15173], wl[15174], wl[15175], wl[15176], wl[15177], wl[15178], wl[15179], wl[15180], wl[15181], wl[15182], wl[15183], wl[15184], wl[15185], wl[15186], wl[15187], wl[15188], wl[15189], wl[15190], wl[15191], wl[15192], wl[15193], wl[15194], wl[15195], wl[15196], wl[15197], wl[15198], wl[15199], wl[15200], wl[15201], wl[15202], wl[15203], wl[15204], wl[15205], wl[15206], wl[15207], wl[15208], wl[15209], wl[15210], wl[15211], wl[15212], wl[15213], wl[15214], wl[15215], wl[15216], wl[15217], wl[15218], wl[15219], wl[15220], wl[15221], wl[15222], wl[15223], wl[17808], wl[17809], wl[17810], wl[17811], wl[17812], wl[17813], wl[17814], wl[17815], wl[17816], wl[17817], wl[17818], wl[17819], wl[17820], wl[17821], wl[17822], wl[17823], wl[17824], wl[17825], wl[17826], wl[17827], wl[17828], wl[17829], wl[17830], wl[17831], wl[17832], wl[17833], wl[17834], wl[17835], wl[17836], wl[17837], wl[17838], wl[17839], wl[17840], wl[17841], wl[17842], wl[17843], wl[17844], wl[17845], wl[17846], wl[17847], wl[17848], wl[17849], wl[17850], wl[17851], wl[17852], wl[17853], wl[17854], wl[17855], wl[17856], wl[17857], wl[17858], wl[17859], wl[17860], wl[17861], wl[17862], wl[17863], wl[17864], wl[17865], wl[17866], wl[17867], wl[17868], wl[17869], wl[17870], wl[17871], wl[17872], wl[17873], wl[17874], wl[17875], wl[17876], wl[17877], wl[17878], wl[17879], wl[17880], wl[17881], wl[17882], wl[17883], wl[17884], wl[17885], wl[17886], wl[17887], wl[14124], wl[14125], wl[14126], wl[14127], wl[14128], wl[14129], wl[14130], wl[14131], wl[14132], wl[14133], wl[14134], wl[14135], wl[14136], wl[14137], wl[14138], wl[14139], wl[14140], wl[14141], wl[14142], wl[14143], wl[14144], wl[14145], wl[14146], wl[14147], wl[14148], wl[14149], wl[14150], wl[14151], wl[14152], wl[14153], wl[14154], wl[14155], wl[14156], wl[14157], wl[14158], wl[14159], wl[14160], wl[14161], wl[14162], wl[14163], wl[14164], wl[14165], wl[14166], wl[14167], wl[14168], wl[14169], wl[14170], wl[14171], wl[14172], wl[14173], wl[14174], wl[14175], wl[14176], wl[14177], wl[14178], wl[14179], wl[14180], wl[14181], wl[14182], wl[14183], wl[14184], wl[14185], wl[14186], wl[14187], wl[14188], wl[14189], wl[14190], wl[14191], wl[14192], wl[14193], wl[14194], wl[14195], wl[14196], wl[14197], wl[14198], wl[14199], wl[14200], wl[14201], wl[14202], wl[14203], wl[17728], wl[17729], wl[17730], wl[17731], wl[17732], wl[17733], wl[17734], wl[17735], wl[17736], wl[17737], wl[17738], wl[17739], wl[17740], wl[17741], wl[17742], wl[17743], wl[17744], wl[17745], wl[17746], wl[17747], wl[17748], wl[17749], wl[17750], wl[17751], wl[17752], wl[17753], wl[17754], wl[17755], wl[17756], wl[17757], wl[17758], wl[17759], wl[17760], wl[17761], wl[17762], wl[17763], wl[17764], wl[17765], wl[17766], wl[17767], wl[17768], wl[17769], wl[17770], wl[17771], wl[17772], wl[17773], wl[17774], wl[17775], wl[17776], wl[17777], wl[17778], wl[17779], wl[17780], wl[17781], wl[17782], wl[17783], wl[17784], wl[17785], wl[17786], wl[17787], wl[17788], wl[17789], wl[17790], wl[17791], wl[17792], wl[17793], wl[17794], wl[17795], wl[17796], wl[17797], wl[17798], wl[17799], wl[17800], wl[17801], wl[17802], wl[17803], wl[17804], wl[17805], wl[17806], wl[17807]})
    );
    right_tile tile_5__2_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_3__1__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_3__1__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_3__1__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_4__0__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_4__0__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_4__0__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_3__0__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_3__0__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_3__0__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_3__0__grid_top_r_in[1]),
        .grid_left_in(grid_clb_4__1__grid_left_in),
        .grid_bottom_in(grid_clb_4__1__grid_bottom_in),
        .chanx_left_in(sb_1__1__6_chanx_right_out),
        .chanx_left_out(cbx_1__1__9_chanx_left_out),
        .grid_top_out(grid_clb_4__2__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[56:63]),
        .io_left_in(grid_io_right_5__1__io_left_in),
        .chany_bottom_in(sb_4__0__0_chany_top_out),
        .chany_bottom_out(cby_4__1__0_chany_bottom_out),
        .chany_top_in_0(cby_4__1__1_chany_bottom_out),
        .chany_top_out_0(sb_4__1__0_chany_top_out),
        .grid_top_r_inpad(grid_io_right_5__2__io_left_in),
        .grid_top_l_in(sb_4__1__grid_top_l_in),
        .grid_bottom_l_in(sb_4__0__grid_top_l_in),
        .grid_left_t_in(sb_3__1__grid_right_t_in),
        .grid_left_b_in(sb_3__1__grid_right_b_in),
        .bl({bl[5392], bl[5393], bl[5394], bl[5395], bl[5396], bl[5397], bl[5398], bl[5399], bl[5400], bl[5401], bl[5402], bl[5403], bl[5404], bl[5405], bl[5406], bl[5407], bl[5408], bl[5409], bl[5410], bl[5411], bl[5412], bl[5413], bl[5414], bl[5415], bl[5416], bl[5417], bl[5418], bl[5419], bl[5420], bl[5421], bl[5422], bl[5423], bl[5424], bl[5425], bl[5426], bl[5427], bl[5428], bl[5429], bl[5430], bl[5431], bl[5432], bl[5433], bl[5434], bl[5435], bl[5436], bl[5437], bl[5438], bl[5439], bl[5440], bl[5441], bl[5442], bl[5443], bl[5444], bl[5445], bl[5446], bl[5447], bl[5448], bl[5449], bl[5450], bl[5451], bl[5452], bl[5453], bl[5454], bl[5455], bl[5456], bl[5457], bl[5458], bl[5459], bl[5460], bl[5461], bl[5462], bl[5463], bl[5464], bl[5465], bl[5466], bl[5467], bl[5468], bl[5469], bl[5470], bl[5471], bl[5472], bl[5473], bl[5474], bl[5475], bl[5476], bl[5477], bl[5478], bl[5479], bl[5480], bl[5481], bl[5482], bl[5483], bl[5484], bl[5485], bl[5486], bl[5487], bl[5488], bl[5489], bl[5490], bl[5491], bl[5492], bl[5493], bl[5494], bl[5495], bl[5496], bl[5497], bl[5498], bl[5499], bl[5500], bl[5501], bl[5502], bl[5503], bl[5504], bl[5505], bl[5506], bl[5507], bl[5508], bl[5509], bl[5510], bl[5511], bl[5512], bl[5513], bl[5514], bl[5515], bl[5516], bl[5517], bl[5518], bl[5519], bl[5520], bl[5521], bl[5522], bl[5523], bl[5524], bl[5525], bl[5526], bl[5527], bl[5528], bl[5529], bl[5530], bl[5531], bl[5532], bl[5533], bl[5534], bl[5535], bl[5536], bl[5537], bl[5538], bl[5539], bl[5540], bl[5541], bl[5542], bl[5543], bl[5544], bl[5545], bl[5546], bl[5547], bl[5548], bl[5549], bl[5550], bl[5551], bl[5552], bl[5553], bl[5554], bl[5555], bl[5556], bl[5557], bl[5558], bl[5559], bl[5560], bl[5561], bl[5562], bl[5563], bl[5564], bl[5565], bl[5566], bl[5567], bl[5568], bl[5569], bl[5570], bl[5571], bl[5572], bl[5573], bl[5574], bl[5575], bl[5576], bl[5577], bl[5578], bl[5579], bl[5580], bl[5581], bl[5582], bl[5583], bl[5584], bl[5585], bl[5586], bl[5587], bl[5588], bl[5589], bl[5590], bl[5591], bl[5592], bl[5593], bl[5594], bl[5595], bl[5596], bl[5597], bl[5598], bl[5599], bl[5600], bl[5601], bl[5602], bl[5603], bl[5604], bl[5605], bl[5606], bl[5607], bl[5608], bl[5609], bl[5610], bl[5611], bl[5612], bl[5613], bl[5614], bl[5615], bl[5616], bl[5617], bl[5618], bl[5619], bl[5620], bl[5621], bl[5622], bl[5623], bl[5624], bl[5625], bl[5626], bl[5627], bl[5628], bl[5629], bl[5630], bl[5631], bl[5632], bl[5633], bl[5634], bl[5635], bl[5636], bl[5637], bl[5638], bl[5639], bl[5640], bl[5641], bl[5642], bl[5643], bl[5644], bl[5645], bl[5646], bl[5647], bl[5648], bl[5649], bl[5650], bl[5651], bl[5652], bl[5653], bl[5654], bl[5655], bl[5656], bl[5657], bl[5658], bl[5659], bl[5660], bl[5661], bl[5662], bl[5663], bl[5664], bl[5665], bl[5666], bl[5667], bl[5668], bl[5669], bl[5670], bl[5671], bl[5672], bl[5673], bl[5674], bl[5675], bl[5676], bl[5677], bl[5678], bl[5679], bl[5680], bl[5681], bl[5682], bl[5683], bl[5684], bl[5685], bl[5686], bl[5687], bl[5688], bl[5689], bl[5690], bl[5691], bl[5692], bl[5693], bl[5694], bl[5695], bl[5696], bl[5697], bl[5698], bl[5699], bl[5700], bl[5701], bl[5702], bl[5703], bl[5704], bl[5705], bl[5706], bl[5707], bl[5708], bl[5709], bl[5710], bl[5711], bl[5712], bl[5713], bl[5714], bl[5715], bl[5716], bl[5717], bl[5718], bl[5719], bl[5720], bl[5721], bl[5722], bl[5723], bl[5724], bl[5725], bl[5726], bl[5727], bl[5728], bl[5729], bl[5730], bl[5731], bl[5732], bl[5733], bl[5734], bl[5735], bl[5736], bl[5737], bl[5738], bl[5739], bl[5740], bl[5741], bl[5742], bl[5743], bl[5744], bl[5745], bl[5746], bl[5747], bl[5748], bl[5749], bl[5750], bl[5751], bl[5752], bl[5753], bl[5754], bl[5755], bl[5756], bl[5757], bl[5758], bl[5759], bl[5760], bl[5761], bl[5762], bl[5763], bl[5764], bl[5765], bl[5766], bl[5767], bl[5768], bl[5769], bl[5770], bl[5771], bl[5772], bl[5773], bl[5774], bl[5775], bl[5776], bl[5777], bl[5778], bl[5779], bl[5780], bl[5781], bl[5782], bl[5783], bl[5784], bl[5785], bl[5786], bl[5787], bl[5788], bl[5789], bl[5790], bl[5791], bl[5792], bl[5793], bl[5794], bl[5795], bl[5796], bl[5797], bl[5798], bl[5799], bl[5800], bl[5801], bl[5802], bl[5803], bl[5804], bl[5805], bl[5806], bl[5807], bl[5808], bl[5809], bl[5810], bl[5811], bl[5812], bl[5813], bl[5814], bl[5815], bl[5816], bl[5817], bl[5818], bl[5819], bl[5820], bl[5821], bl[5822], bl[5823], bl[5824], bl[5825], bl[5826], bl[5827], bl[5828], bl[5829], bl[5830], bl[5831], bl[5832], bl[5833], bl[5834], bl[5835], bl[5836], bl[5837], bl[5838], bl[5839], bl[5840], bl[5841], bl[5842], bl[5843], bl[5844], bl[5845], bl[5846], bl[5847], bl[5848], bl[5849], bl[5850], bl[5851], bl[5852], bl[5853], bl[5854], bl[5855], bl[5856], bl[5857], bl[5858], bl[5859], bl[5860], bl[5861], bl[5862], bl[5863], bl[5864], bl[5865], bl[5866], bl[5867], bl[5868], bl[5869], bl[5870], bl[5871], bl[5872], bl[5873], bl[5874], bl[5875], bl[5876], bl[5877], bl[5878], bl[5879], bl[5880], bl[5881], bl[5882], bl[5883], bl[5884], bl[5885], bl[5886], bl[5887], bl[5888], bl[5889], bl[5890], bl[5891], bl[5892], bl[5893], bl[5894], bl[5895], bl[5896], bl[5897], bl[5898], bl[5899], bl[5900], bl[5901], bl[5902], bl[5903], bl[5904], bl[5905], bl[5906], bl[5907], bl[5908], bl[5909], bl[5910], bl[5911], bl[5912], bl[5913], bl[5914], bl[5915], bl[5916], bl[5917], bl[5918], bl[5919], bl[5920], bl[5921], bl[5922], bl[5923], bl[5924], bl[5925], bl[5926], bl[5927], bl[5928], bl[5929], bl[5930], bl[5931], bl[5932], bl[5933], bl[5934], bl[5935], bl[5936], bl[5937], bl[5938], bl[5939], bl[5940], bl[5941], bl[5942], bl[5943], bl[5944], bl[5945], bl[5946], bl[5947], bl[5948], bl[5949], bl[5950], bl[5951], bl[5952], bl[5953], bl[5954], bl[5955], bl[5956], bl[5957], bl[5958], bl[5959], bl[5960], bl[5961], bl[5962], bl[5963], bl[5964], bl[5965], bl[5966], bl[5967], bl[5968], bl[5969], bl[5970], bl[5971], bl[5972], bl[5973], bl[5974], bl[5975], bl[5976], bl[5977], bl[5978], bl[5979], bl[5980], bl[5981], bl[5982], bl[5983], bl[5984], bl[5985], bl[5986], bl[5987], bl[5988], bl[5989], bl[5990], bl[5991], bl[5992], bl[5993], bl[5994], bl[5995], bl[5996], bl[5997], bl[5998], bl[5999], bl[6000], bl[6001], bl[6002], bl[6003], bl[6004], bl[6005], bl[6006], bl[6007], bl[6008], bl[6009], bl[6010], bl[6011], bl[6012], bl[6013], bl[6014], bl[6015], bl[6016], bl[6017], bl[6018], bl[6019], bl[6020], bl[6021], bl[6022], bl[6023], bl[6024], bl[6025], bl[6026], bl[6027], bl[6028], bl[6029], bl[6030], bl[6031], bl[6032], bl[6033], bl[6034], bl[6035], bl[6036], bl[6037], bl[6038], bl[6039], bl[6040], bl[6041], bl[6042], bl[6043], bl[6044], bl[6045], bl[6046], bl[6047], bl[6048], bl[6049], bl[6050], bl[6051], bl[6052], bl[6053], bl[6054], bl[6055], bl[6056], bl[6057], bl[6058], bl[6059], bl[6060], bl[6061], bl[6062], bl[6063], bl[6064], bl[6065], bl[6066], bl[6067], bl[6068], bl[6069], bl[6070], bl[6071], bl[6072], bl[6073], bl[6074], bl[6075], bl[6076], bl[6077], bl[6078], bl[6079], bl[6080], bl[6081], bl[6082], bl[6083], bl[6084], bl[6085], bl[6086], bl[6087], bl[6088], bl[6089], bl[6090], bl[6091], bl[6092], bl[6093], bl[6094], bl[6095], bl[6096], bl[6097], bl[6098], bl[6099], bl[6100], bl[6101], bl[6102], bl[6103], bl[6104], bl[6105], bl[6106], bl[6107], bl[6108], bl[6109], bl[6110], bl[6111], bl[6112], bl[6113], bl[6114], bl[6115], bl[6116], bl[6117], bl[6118], bl[6119], bl[6120], bl[6121], bl[6122], bl[6123], bl[6124], bl[6125], bl[6126], bl[6127], bl[6128], bl[6129], bl[6130], bl[6131], bl[6132], bl[6133], bl[6134], bl[6135], bl[6136], bl[6137], bl[6138], bl[6139], bl[6140], bl[6141], bl[6142], bl[6143], bl[6144], bl[6145], bl[6146], bl[6147], bl[6148], bl[6149], bl[6150], bl[6151], bl[6152], bl[6153], bl[6154], bl[6155], bl[6156], bl[6157], bl[6158], bl[6159], bl[6160], bl[6161], bl[6162], bl[6163], bl[6164], bl[6165], bl[6166], bl[6167], bl[6168], bl[6169], bl[6170], bl[6171], bl[6172], bl[6173], bl[6174], bl[6175], bl[6176], bl[6177], bl[6178], bl[6179], bl[6180], bl[6181], bl[6182], bl[6183], bl[6184], bl[6185], bl[6186], bl[6187], bl[6188], bl[6189], bl[6190], bl[6191], bl[6192], bl[6193], bl[6194], bl[6195], bl[6196], bl[6197], bl[6198], bl[6199], bl[6200], bl[6201], bl[6202], bl[6203], bl[6204], bl[6205], bl[6206], bl[6207], bl[6208], bl[6209], bl[6210], bl[6211], bl[6212], bl[6213], bl[6214], bl[6215], bl[6216], bl[6217], bl[6218], bl[6219], bl[6220], bl[6221], bl[6222], bl[6223], bl[6224], bl[6225], bl[6226], bl[6227], bl[6228], bl[6229], bl[6230], bl[6231], bl[6232], bl[6233], bl[6234], bl[6235], bl[6236], bl[6237], bl[6238], bl[6239], bl[6240], bl[6241], bl[6242], bl[6243], bl[6244], bl[6245], bl[6246], bl[6247], bl[6248], bl[6249], bl[6250], bl[6251], bl[6252], bl[6253], bl[6254], bl[6255], bl[6256], bl[6257], bl[6258], bl[6259], bl[6260], bl[6261], bl[6262], bl[6263], bl[6264], bl[6265], bl[6266], bl[6267], bl[6268], bl[6269], bl[6270], bl[6271], bl[6272], bl[6273], bl[6274], bl[6275], bl[6276], bl[6277], bl[6278], bl[6279], bl[6280], bl[6281], bl[6282], bl[6283], bl[6284], bl[6285], bl[6286], bl[6287], bl[6288], bl[6289], bl[6290], bl[6291], bl[6292], bl[6293], bl[6294], bl[6295], bl[6296], bl[6297], bl[6298], bl[6299], bl[6300], bl[6301], bl[6302], bl[6303], bl[6304], bl[6305], bl[6306], bl[6307], bl[6308], bl[6309], bl[6310], bl[6311], bl[6312], bl[6313], bl[6314], bl[6315], bl[6316], bl[6317], bl[6318], bl[6319], bl[6320], bl[6321], bl[6322], bl[6323], bl[6324], bl[6325], bl[6326], bl[6327], bl[6328], bl[6329], bl[6330], bl[6331], bl[6332], bl[6333], bl[6334], bl[6335], bl[6336], bl[6337], bl[6338], bl[6339], bl[6340], bl[6341], bl[6342], bl[6343], bl[6344], bl[6345], bl[6346], bl[6347], bl[6348], bl[6349], bl[6350], bl[6351], bl[6352], bl[6353], bl[6354], bl[6355], bl[6356], bl[6357], bl[6358], bl[6359], bl[6360], bl[6361], bl[6362], bl[6363], bl[6364], bl[6365], bl[6366], bl[6367], bl[6368], bl[6369], bl[6370], bl[6371], bl[6372], bl[6373], bl[6374], bl[6375], bl[6376], bl[6377], bl[6378], bl[6379], bl[6380], bl[6381], bl[6382], bl[6383], bl[6384], bl[6385], bl[6386], bl[6387], bl[6388], bl[6389], bl[6390], bl[6391], bl[6392], bl[6393], bl[6394], bl[6395], bl[6396], bl[6397], bl[6398], bl[6399], bl[6400], bl[6401], bl[6402], bl[6403], bl[6404], bl[6405], bl[6406], bl[6407], bl[6408], bl[6409], bl[6410], bl[6411], bl[6492], bl[6493], bl[6494], bl[6495], bl[6496], bl[6497], bl[6498], bl[6499], bl[6500], bl[6501], bl[6502], bl[6503], bl[6504], bl[6505], bl[6506], bl[6507], bl[6508], bl[6509], bl[6510], bl[6511], bl[6512], bl[6513], bl[6514], bl[6515], bl[6516], bl[6517], bl[6518], bl[6519], bl[6520], bl[6521], bl[6522], bl[6523], bl[6524], bl[6525], bl[6526], bl[6527], bl[6528], bl[6529], bl[6530], bl[6531], bl[6532], bl[6533], bl[6534], bl[6535], bl[6536], bl[6537], bl[6538], bl[6539], bl[6540], bl[6541], bl[6542], bl[6543], bl[6544], bl[6545], bl[6546], bl[6547], bl[6548], bl[6549], bl[6550], bl[6551], bl[6552], bl[6553], bl[6554], bl[6555], bl[6556], bl[6557], bl[6558], bl[6559], bl[6560], bl[6561], bl[6562], bl[6563], bl[6564], bl[6565], bl[6566], bl[6567], bl[6568], bl[6569], bl[6570], bl[6571], bl[32], bl[33], bl[34], bl[35], bl[36], bl[37], bl[38], bl[39], bl[5320], bl[5321], bl[5322], bl[5323], bl[5324], bl[5325], bl[5326], bl[5327], bl[5328], bl[5329], bl[5330], bl[5331], bl[5332], bl[5333], bl[5334], bl[5335], bl[5336], bl[5337], bl[5338], bl[5339], bl[5340], bl[5341], bl[5342], bl[5343], bl[5344], bl[5345], bl[5346], bl[5347], bl[5348], bl[5349], bl[5350], bl[5351], bl[5352], bl[5353], bl[5354], bl[5355], bl[5356], bl[5357], bl[5358], bl[5359], bl[5360], bl[5361], bl[5362], bl[5363], bl[5364], bl[5365], bl[5366], bl[5367], bl[5368], bl[5369], bl[5370], bl[5371], bl[5372], bl[5373], bl[5374], bl[5375], bl[5376], bl[5377], bl[5378], bl[5379], bl[5380], bl[5381], bl[5382], bl[5383], bl[5384], bl[5385], bl[5386], bl[5387], bl[5388], bl[5389], bl[5390], bl[5391], bl[6412], bl[6413], bl[6414], bl[6415], bl[6416], bl[6417], bl[6418], bl[6419], bl[6420], bl[6421], bl[6422], bl[6423], bl[6424], bl[6425], bl[6426], bl[6427], bl[6428], bl[6429], bl[6430], bl[6431], bl[6432], bl[6433], bl[6434], bl[6435], bl[6436], bl[6437], bl[6438], bl[6439], bl[6440], bl[6441], bl[6442], bl[6443], bl[6444], bl[6445], bl[6446], bl[6447], bl[6448], bl[6449], bl[6450], bl[6451], bl[6452], bl[6453], bl[6454], bl[6455], bl[6456], bl[6457], bl[6458], bl[6459], bl[6460], bl[6461], bl[6462], bl[6463], bl[6464], bl[6465], bl[6466], bl[6467], bl[6468], bl[6469], bl[6470], bl[6471], bl[6472], bl[6473], bl[6474], bl[6475], bl[6476], bl[6477], bl[6478], bl[6479], bl[6480], bl[6481], bl[6482], bl[6483], bl[6484], bl[6485], bl[6486], bl[6487], bl[6488], bl[6489], bl[6490], bl[6491]}),
        .wl({wl[5392], wl[5393], wl[5394], wl[5395], wl[5396], wl[5397], wl[5398], wl[5399], wl[5400], wl[5401], wl[5402], wl[5403], wl[5404], wl[5405], wl[5406], wl[5407], wl[5408], wl[5409], wl[5410], wl[5411], wl[5412], wl[5413], wl[5414], wl[5415], wl[5416], wl[5417], wl[5418], wl[5419], wl[5420], wl[5421], wl[5422], wl[5423], wl[5424], wl[5425], wl[5426], wl[5427], wl[5428], wl[5429], wl[5430], wl[5431], wl[5432], wl[5433], wl[5434], wl[5435], wl[5436], wl[5437], wl[5438], wl[5439], wl[5440], wl[5441], wl[5442], wl[5443], wl[5444], wl[5445], wl[5446], wl[5447], wl[5448], wl[5449], wl[5450], wl[5451], wl[5452], wl[5453], wl[5454], wl[5455], wl[5456], wl[5457], wl[5458], wl[5459], wl[5460], wl[5461], wl[5462], wl[5463], wl[5464], wl[5465], wl[5466], wl[5467], wl[5468], wl[5469], wl[5470], wl[5471], wl[5472], wl[5473], wl[5474], wl[5475], wl[5476], wl[5477], wl[5478], wl[5479], wl[5480], wl[5481], wl[5482], wl[5483], wl[5484], wl[5485], wl[5486], wl[5487], wl[5488], wl[5489], wl[5490], wl[5491], wl[5492], wl[5493], wl[5494], wl[5495], wl[5496], wl[5497], wl[5498], wl[5499], wl[5500], wl[5501], wl[5502], wl[5503], wl[5504], wl[5505], wl[5506], wl[5507], wl[5508], wl[5509], wl[5510], wl[5511], wl[5512], wl[5513], wl[5514], wl[5515], wl[5516], wl[5517], wl[5518], wl[5519], wl[5520], wl[5521], wl[5522], wl[5523], wl[5524], wl[5525], wl[5526], wl[5527], wl[5528], wl[5529], wl[5530], wl[5531], wl[5532], wl[5533], wl[5534], wl[5535], wl[5536], wl[5537], wl[5538], wl[5539], wl[5540], wl[5541], wl[5542], wl[5543], wl[5544], wl[5545], wl[5546], wl[5547], wl[5548], wl[5549], wl[5550], wl[5551], wl[5552], wl[5553], wl[5554], wl[5555], wl[5556], wl[5557], wl[5558], wl[5559], wl[5560], wl[5561], wl[5562], wl[5563], wl[5564], wl[5565], wl[5566], wl[5567], wl[5568], wl[5569], wl[5570], wl[5571], wl[5572], wl[5573], wl[5574], wl[5575], wl[5576], wl[5577], wl[5578], wl[5579], wl[5580], wl[5581], wl[5582], wl[5583], wl[5584], wl[5585], wl[5586], wl[5587], wl[5588], wl[5589], wl[5590], wl[5591], wl[5592], wl[5593], wl[5594], wl[5595], wl[5596], wl[5597], wl[5598], wl[5599], wl[5600], wl[5601], wl[5602], wl[5603], wl[5604], wl[5605], wl[5606], wl[5607], wl[5608], wl[5609], wl[5610], wl[5611], wl[5612], wl[5613], wl[5614], wl[5615], wl[5616], wl[5617], wl[5618], wl[5619], wl[5620], wl[5621], wl[5622], wl[5623], wl[5624], wl[5625], wl[5626], wl[5627], wl[5628], wl[5629], wl[5630], wl[5631], wl[5632], wl[5633], wl[5634], wl[5635], wl[5636], wl[5637], wl[5638], wl[5639], wl[5640], wl[5641], wl[5642], wl[5643], wl[5644], wl[5645], wl[5646], wl[5647], wl[5648], wl[5649], wl[5650], wl[5651], wl[5652], wl[5653], wl[5654], wl[5655], wl[5656], wl[5657], wl[5658], wl[5659], wl[5660], wl[5661], wl[5662], wl[5663], wl[5664], wl[5665], wl[5666], wl[5667], wl[5668], wl[5669], wl[5670], wl[5671], wl[5672], wl[5673], wl[5674], wl[5675], wl[5676], wl[5677], wl[5678], wl[5679], wl[5680], wl[5681], wl[5682], wl[5683], wl[5684], wl[5685], wl[5686], wl[5687], wl[5688], wl[5689], wl[5690], wl[5691], wl[5692], wl[5693], wl[5694], wl[5695], wl[5696], wl[5697], wl[5698], wl[5699], wl[5700], wl[5701], wl[5702], wl[5703], wl[5704], wl[5705], wl[5706], wl[5707], wl[5708], wl[5709], wl[5710], wl[5711], wl[5712], wl[5713], wl[5714], wl[5715], wl[5716], wl[5717], wl[5718], wl[5719], wl[5720], wl[5721], wl[5722], wl[5723], wl[5724], wl[5725], wl[5726], wl[5727], wl[5728], wl[5729], wl[5730], wl[5731], wl[5732], wl[5733], wl[5734], wl[5735], wl[5736], wl[5737], wl[5738], wl[5739], wl[5740], wl[5741], wl[5742], wl[5743], wl[5744], wl[5745], wl[5746], wl[5747], wl[5748], wl[5749], wl[5750], wl[5751], wl[5752], wl[5753], wl[5754], wl[5755], wl[5756], wl[5757], wl[5758], wl[5759], wl[5760], wl[5761], wl[5762], wl[5763], wl[5764], wl[5765], wl[5766], wl[5767], wl[5768], wl[5769], wl[5770], wl[5771], wl[5772], wl[5773], wl[5774], wl[5775], wl[5776], wl[5777], wl[5778], wl[5779], wl[5780], wl[5781], wl[5782], wl[5783], wl[5784], wl[5785], wl[5786], wl[5787], wl[5788], wl[5789], wl[5790], wl[5791], wl[5792], wl[5793], wl[5794], wl[5795], wl[5796], wl[5797], wl[5798], wl[5799], wl[5800], wl[5801], wl[5802], wl[5803], wl[5804], wl[5805], wl[5806], wl[5807], wl[5808], wl[5809], wl[5810], wl[5811], wl[5812], wl[5813], wl[5814], wl[5815], wl[5816], wl[5817], wl[5818], wl[5819], wl[5820], wl[5821], wl[5822], wl[5823], wl[5824], wl[5825], wl[5826], wl[5827], wl[5828], wl[5829], wl[5830], wl[5831], wl[5832], wl[5833], wl[5834], wl[5835], wl[5836], wl[5837], wl[5838], wl[5839], wl[5840], wl[5841], wl[5842], wl[5843], wl[5844], wl[5845], wl[5846], wl[5847], wl[5848], wl[5849], wl[5850], wl[5851], wl[5852], wl[5853], wl[5854], wl[5855], wl[5856], wl[5857], wl[5858], wl[5859], wl[5860], wl[5861], wl[5862], wl[5863], wl[5864], wl[5865], wl[5866], wl[5867], wl[5868], wl[5869], wl[5870], wl[5871], wl[5872], wl[5873], wl[5874], wl[5875], wl[5876], wl[5877], wl[5878], wl[5879], wl[5880], wl[5881], wl[5882], wl[5883], wl[5884], wl[5885], wl[5886], wl[5887], wl[5888], wl[5889], wl[5890], wl[5891], wl[5892], wl[5893], wl[5894], wl[5895], wl[5896], wl[5897], wl[5898], wl[5899], wl[5900], wl[5901], wl[5902], wl[5903], wl[5904], wl[5905], wl[5906], wl[5907], wl[5908], wl[5909], wl[5910], wl[5911], wl[5912], wl[5913], wl[5914], wl[5915], wl[5916], wl[5917], wl[5918], wl[5919], wl[5920], wl[5921], wl[5922], wl[5923], wl[5924], wl[5925], wl[5926], wl[5927], wl[5928], wl[5929], wl[5930], wl[5931], wl[5932], wl[5933], wl[5934], wl[5935], wl[5936], wl[5937], wl[5938], wl[5939], wl[5940], wl[5941], wl[5942], wl[5943], wl[5944], wl[5945], wl[5946], wl[5947], wl[5948], wl[5949], wl[5950], wl[5951], wl[5952], wl[5953], wl[5954], wl[5955], wl[5956], wl[5957], wl[5958], wl[5959], wl[5960], wl[5961], wl[5962], wl[5963], wl[5964], wl[5965], wl[5966], wl[5967], wl[5968], wl[5969], wl[5970], wl[5971], wl[5972], wl[5973], wl[5974], wl[5975], wl[5976], wl[5977], wl[5978], wl[5979], wl[5980], wl[5981], wl[5982], wl[5983], wl[5984], wl[5985], wl[5986], wl[5987], wl[5988], wl[5989], wl[5990], wl[5991], wl[5992], wl[5993], wl[5994], wl[5995], wl[5996], wl[5997], wl[5998], wl[5999], wl[6000], wl[6001], wl[6002], wl[6003], wl[6004], wl[6005], wl[6006], wl[6007], wl[6008], wl[6009], wl[6010], wl[6011], wl[6012], wl[6013], wl[6014], wl[6015], wl[6016], wl[6017], wl[6018], wl[6019], wl[6020], wl[6021], wl[6022], wl[6023], wl[6024], wl[6025], wl[6026], wl[6027], wl[6028], wl[6029], wl[6030], wl[6031], wl[6032], wl[6033], wl[6034], wl[6035], wl[6036], wl[6037], wl[6038], wl[6039], wl[6040], wl[6041], wl[6042], wl[6043], wl[6044], wl[6045], wl[6046], wl[6047], wl[6048], wl[6049], wl[6050], wl[6051], wl[6052], wl[6053], wl[6054], wl[6055], wl[6056], wl[6057], wl[6058], wl[6059], wl[6060], wl[6061], wl[6062], wl[6063], wl[6064], wl[6065], wl[6066], wl[6067], wl[6068], wl[6069], wl[6070], wl[6071], wl[6072], wl[6073], wl[6074], wl[6075], wl[6076], wl[6077], wl[6078], wl[6079], wl[6080], wl[6081], wl[6082], wl[6083], wl[6084], wl[6085], wl[6086], wl[6087], wl[6088], wl[6089], wl[6090], wl[6091], wl[6092], wl[6093], wl[6094], wl[6095], wl[6096], wl[6097], wl[6098], wl[6099], wl[6100], wl[6101], wl[6102], wl[6103], wl[6104], wl[6105], wl[6106], wl[6107], wl[6108], wl[6109], wl[6110], wl[6111], wl[6112], wl[6113], wl[6114], wl[6115], wl[6116], wl[6117], wl[6118], wl[6119], wl[6120], wl[6121], wl[6122], wl[6123], wl[6124], wl[6125], wl[6126], wl[6127], wl[6128], wl[6129], wl[6130], wl[6131], wl[6132], wl[6133], wl[6134], wl[6135], wl[6136], wl[6137], wl[6138], wl[6139], wl[6140], wl[6141], wl[6142], wl[6143], wl[6144], wl[6145], wl[6146], wl[6147], wl[6148], wl[6149], wl[6150], wl[6151], wl[6152], wl[6153], wl[6154], wl[6155], wl[6156], wl[6157], wl[6158], wl[6159], wl[6160], wl[6161], wl[6162], wl[6163], wl[6164], wl[6165], wl[6166], wl[6167], wl[6168], wl[6169], wl[6170], wl[6171], wl[6172], wl[6173], wl[6174], wl[6175], wl[6176], wl[6177], wl[6178], wl[6179], wl[6180], wl[6181], wl[6182], wl[6183], wl[6184], wl[6185], wl[6186], wl[6187], wl[6188], wl[6189], wl[6190], wl[6191], wl[6192], wl[6193], wl[6194], wl[6195], wl[6196], wl[6197], wl[6198], wl[6199], wl[6200], wl[6201], wl[6202], wl[6203], wl[6204], wl[6205], wl[6206], wl[6207], wl[6208], wl[6209], wl[6210], wl[6211], wl[6212], wl[6213], wl[6214], wl[6215], wl[6216], wl[6217], wl[6218], wl[6219], wl[6220], wl[6221], wl[6222], wl[6223], wl[6224], wl[6225], wl[6226], wl[6227], wl[6228], wl[6229], wl[6230], wl[6231], wl[6232], wl[6233], wl[6234], wl[6235], wl[6236], wl[6237], wl[6238], wl[6239], wl[6240], wl[6241], wl[6242], wl[6243], wl[6244], wl[6245], wl[6246], wl[6247], wl[6248], wl[6249], wl[6250], wl[6251], wl[6252], wl[6253], wl[6254], wl[6255], wl[6256], wl[6257], wl[6258], wl[6259], wl[6260], wl[6261], wl[6262], wl[6263], wl[6264], wl[6265], wl[6266], wl[6267], wl[6268], wl[6269], wl[6270], wl[6271], wl[6272], wl[6273], wl[6274], wl[6275], wl[6276], wl[6277], wl[6278], wl[6279], wl[6280], wl[6281], wl[6282], wl[6283], wl[6284], wl[6285], wl[6286], wl[6287], wl[6288], wl[6289], wl[6290], wl[6291], wl[6292], wl[6293], wl[6294], wl[6295], wl[6296], wl[6297], wl[6298], wl[6299], wl[6300], wl[6301], wl[6302], wl[6303], wl[6304], wl[6305], wl[6306], wl[6307], wl[6308], wl[6309], wl[6310], wl[6311], wl[6312], wl[6313], wl[6314], wl[6315], wl[6316], wl[6317], wl[6318], wl[6319], wl[6320], wl[6321], wl[6322], wl[6323], wl[6324], wl[6325], wl[6326], wl[6327], wl[6328], wl[6329], wl[6330], wl[6331], wl[6332], wl[6333], wl[6334], wl[6335], wl[6336], wl[6337], wl[6338], wl[6339], wl[6340], wl[6341], wl[6342], wl[6343], wl[6344], wl[6345], wl[6346], wl[6347], wl[6348], wl[6349], wl[6350], wl[6351], wl[6352], wl[6353], wl[6354], wl[6355], wl[6356], wl[6357], wl[6358], wl[6359], wl[6360], wl[6361], wl[6362], wl[6363], wl[6364], wl[6365], wl[6366], wl[6367], wl[6368], wl[6369], wl[6370], wl[6371], wl[6372], wl[6373], wl[6374], wl[6375], wl[6376], wl[6377], wl[6378], wl[6379], wl[6380], wl[6381], wl[6382], wl[6383], wl[6384], wl[6385], wl[6386], wl[6387], wl[6388], wl[6389], wl[6390], wl[6391], wl[6392], wl[6393], wl[6394], wl[6395], wl[6396], wl[6397], wl[6398], wl[6399], wl[6400], wl[6401], wl[6402], wl[6403], wl[6404], wl[6405], wl[6406], wl[6407], wl[6408], wl[6409], wl[6410], wl[6411], wl[6492], wl[6493], wl[6494], wl[6495], wl[6496], wl[6497], wl[6498], wl[6499], wl[6500], wl[6501], wl[6502], wl[6503], wl[6504], wl[6505], wl[6506], wl[6507], wl[6508], wl[6509], wl[6510], wl[6511], wl[6512], wl[6513], wl[6514], wl[6515], wl[6516], wl[6517], wl[6518], wl[6519], wl[6520], wl[6521], wl[6522], wl[6523], wl[6524], wl[6525], wl[6526], wl[6527], wl[6528], wl[6529], wl[6530], wl[6531], wl[6532], wl[6533], wl[6534], wl[6535], wl[6536], wl[6537], wl[6538], wl[6539], wl[6540], wl[6541], wl[6542], wl[6543], wl[6544], wl[6545], wl[6546], wl[6547], wl[6548], wl[6549], wl[6550], wl[6551], wl[6552], wl[6553], wl[6554], wl[6555], wl[6556], wl[6557], wl[6558], wl[6559], wl[6560], wl[6561], wl[6562], wl[6563], wl[6564], wl[6565], wl[6566], wl[6567], wl[6568], wl[6569], wl[6570], wl[6571], wl[32], wl[33], wl[34], wl[35], wl[36], wl[37], wl[38], wl[39], wl[5320], wl[5321], wl[5322], wl[5323], wl[5324], wl[5325], wl[5326], wl[5327], wl[5328], wl[5329], wl[5330], wl[5331], wl[5332], wl[5333], wl[5334], wl[5335], wl[5336], wl[5337], wl[5338], wl[5339], wl[5340], wl[5341], wl[5342], wl[5343], wl[5344], wl[5345], wl[5346], wl[5347], wl[5348], wl[5349], wl[5350], wl[5351], wl[5352], wl[5353], wl[5354], wl[5355], wl[5356], wl[5357], wl[5358], wl[5359], wl[5360], wl[5361], wl[5362], wl[5363], wl[5364], wl[5365], wl[5366], wl[5367], wl[5368], wl[5369], wl[5370], wl[5371], wl[5372], wl[5373], wl[5374], wl[5375], wl[5376], wl[5377], wl[5378], wl[5379], wl[5380], wl[5381], wl[5382], wl[5383], wl[5384], wl[5385], wl[5386], wl[5387], wl[5388], wl[5389], wl[5390], wl[5391], wl[6412], wl[6413], wl[6414], wl[6415], wl[6416], wl[6417], wl[6418], wl[6419], wl[6420], wl[6421], wl[6422], wl[6423], wl[6424], wl[6425], wl[6426], wl[6427], wl[6428], wl[6429], wl[6430], wl[6431], wl[6432], wl[6433], wl[6434], wl[6435], wl[6436], wl[6437], wl[6438], wl[6439], wl[6440], wl[6441], wl[6442], wl[6443], wl[6444], wl[6445], wl[6446], wl[6447], wl[6448], wl[6449], wl[6450], wl[6451], wl[6452], wl[6453], wl[6454], wl[6455], wl[6456], wl[6457], wl[6458], wl[6459], wl[6460], wl[6461], wl[6462], wl[6463], wl[6464], wl[6465], wl[6466], wl[6467], wl[6468], wl[6469], wl[6470], wl[6471], wl[6472], wl[6473], wl[6474], wl[6475], wl[6476], wl[6477], wl[6478], wl[6479], wl[6480], wl[6481], wl[6482], wl[6483], wl[6484], wl[6485], wl[6486], wl[6487], wl[6488], wl[6489], wl[6490], wl[6491]})
    );
    right_tile tile_5__3_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_3__2__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_3__2__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_3__2__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_4__1__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_4__1__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_4__1__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_3__1__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_3__1__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_3__1__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_3__1__grid_top_r_in[1]),
        .grid_left_in(grid_clb_4__2__grid_left_in),
        .grid_bottom_in(grid_clb_4__2__grid_bottom_in),
        .chanx_left_in(sb_1__1__7_chanx_right_out),
        .chanx_left_out(cbx_1__1__10_chanx_left_out),
        .grid_top_out(grid_clb_4__3__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[48:55]),
        .io_left_in(grid_io_right_5__2__io_left_in),
        .chany_bottom_in(sb_4__1__0_chany_top_out),
        .chany_bottom_out(cby_4__1__1_chany_bottom_out),
        .chany_top_in_0(cby_4__1__2_chany_bottom_out),
        .chany_top_out_0(sb_4__1__1_chany_top_out),
        .grid_top_r_inpad(grid_io_right_5__3__io_left_in),
        .grid_top_l_in(sb_4__2__grid_top_l_in),
        .grid_bottom_l_in(sb_4__1__grid_top_l_in),
        .grid_left_t_in(sb_3__2__grid_right_t_in),
        .grid_left_b_in(sb_3__2__grid_right_b_in),
        .bl({bl[6644], bl[6645], bl[6646], bl[6647], bl[6648], bl[6649], bl[6650], bl[6651], bl[6652], bl[6653], bl[6654], bl[6655], bl[6656], bl[6657], bl[6658], bl[6659], bl[6660], bl[6661], bl[6662], bl[6663], bl[6664], bl[6665], bl[6666], bl[6667], bl[6668], bl[6669], bl[6670], bl[6671], bl[6672], bl[6673], bl[6674], bl[6675], bl[6676], bl[6677], bl[6678], bl[6679], bl[6680], bl[6681], bl[6682], bl[6683], bl[6684], bl[6685], bl[6686], bl[6687], bl[6688], bl[6689], bl[6690], bl[6691], bl[6692], bl[6693], bl[6694], bl[6695], bl[6696], bl[6697], bl[6698], bl[6699], bl[6700], bl[6701], bl[6702], bl[6703], bl[6704], bl[6705], bl[6706], bl[6707], bl[6708], bl[6709], bl[6710], bl[6711], bl[6712], bl[6713], bl[6714], bl[6715], bl[6716], bl[6717], bl[6718], bl[6719], bl[6720], bl[6721], bl[6722], bl[6723], bl[6724], bl[6725], bl[6726], bl[6727], bl[6728], bl[6729], bl[6730], bl[6731], bl[6732], bl[6733], bl[6734], bl[6735], bl[6736], bl[6737], bl[6738], bl[6739], bl[6740], bl[6741], bl[6742], bl[6743], bl[6744], bl[6745], bl[6746], bl[6747], bl[6748], bl[6749], bl[6750], bl[6751], bl[6752], bl[6753], bl[6754], bl[6755], bl[6756], bl[6757], bl[6758], bl[6759], bl[6760], bl[6761], bl[6762], bl[6763], bl[6764], bl[6765], bl[6766], bl[6767], bl[6768], bl[6769], bl[6770], bl[6771], bl[6772], bl[6773], bl[6774], bl[6775], bl[6776], bl[6777], bl[6778], bl[6779], bl[6780], bl[6781], bl[6782], bl[6783], bl[6784], bl[6785], bl[6786], bl[6787], bl[6788], bl[6789], bl[6790], bl[6791], bl[6792], bl[6793], bl[6794], bl[6795], bl[6796], bl[6797], bl[6798], bl[6799], bl[6800], bl[6801], bl[6802], bl[6803], bl[6804], bl[6805], bl[6806], bl[6807], bl[6808], bl[6809], bl[6810], bl[6811], bl[6812], bl[6813], bl[6814], bl[6815], bl[6816], bl[6817], bl[6818], bl[6819], bl[6820], bl[6821], bl[6822], bl[6823], bl[6824], bl[6825], bl[6826], bl[6827], bl[6828], bl[6829], bl[6830], bl[6831], bl[6832], bl[6833], bl[6834], bl[6835], bl[6836], bl[6837], bl[6838], bl[6839], bl[6840], bl[6841], bl[6842], bl[6843], bl[6844], bl[6845], bl[6846], bl[6847], bl[6848], bl[6849], bl[6850], bl[6851], bl[6852], bl[6853], bl[6854], bl[6855], bl[6856], bl[6857], bl[6858], bl[6859], bl[6860], bl[6861], bl[6862], bl[6863], bl[6864], bl[6865], bl[6866], bl[6867], bl[6868], bl[6869], bl[6870], bl[6871], bl[6872], bl[6873], bl[6874], bl[6875], bl[6876], bl[6877], bl[6878], bl[6879], bl[6880], bl[6881], bl[6882], bl[6883], bl[6884], bl[6885], bl[6886], bl[6887], bl[6888], bl[6889], bl[6890], bl[6891], bl[6892], bl[6893], bl[6894], bl[6895], bl[6896], bl[6897], bl[6898], bl[6899], bl[6900], bl[6901], bl[6902], bl[6903], bl[6904], bl[6905], bl[6906], bl[6907], bl[6908], bl[6909], bl[6910], bl[6911], bl[6912], bl[6913], bl[6914], bl[6915], bl[6916], bl[6917], bl[6918], bl[6919], bl[6920], bl[6921], bl[6922], bl[6923], bl[6924], bl[6925], bl[6926], bl[6927], bl[6928], bl[6929], bl[6930], bl[6931], bl[6932], bl[6933], bl[6934], bl[6935], bl[6936], bl[6937], bl[6938], bl[6939], bl[6940], bl[6941], bl[6942], bl[6943], bl[6944], bl[6945], bl[6946], bl[6947], bl[6948], bl[6949], bl[6950], bl[6951], bl[6952], bl[6953], bl[6954], bl[6955], bl[6956], bl[6957], bl[6958], bl[6959], bl[6960], bl[6961], bl[6962], bl[6963], bl[6964], bl[6965], bl[6966], bl[6967], bl[6968], bl[6969], bl[6970], bl[6971], bl[6972], bl[6973], bl[6974], bl[6975], bl[6976], bl[6977], bl[6978], bl[6979], bl[6980], bl[6981], bl[6982], bl[6983], bl[6984], bl[6985], bl[6986], bl[6987], bl[6988], bl[6989], bl[6990], bl[6991], bl[6992], bl[6993], bl[6994], bl[6995], bl[6996], bl[6997], bl[6998], bl[6999], bl[7000], bl[7001], bl[7002], bl[7003], bl[7004], bl[7005], bl[7006], bl[7007], bl[7008], bl[7009], bl[7010], bl[7011], bl[7012], bl[7013], bl[7014], bl[7015], bl[7016], bl[7017], bl[7018], bl[7019], bl[7020], bl[7021], bl[7022], bl[7023], bl[7024], bl[7025], bl[7026], bl[7027], bl[7028], bl[7029], bl[7030], bl[7031], bl[7032], bl[7033], bl[7034], bl[7035], bl[7036], bl[7037], bl[7038], bl[7039], bl[7040], bl[7041], bl[7042], bl[7043], bl[7044], bl[7045], bl[7046], bl[7047], bl[7048], bl[7049], bl[7050], bl[7051], bl[7052], bl[7053], bl[7054], bl[7055], bl[7056], bl[7057], bl[7058], bl[7059], bl[7060], bl[7061], bl[7062], bl[7063], bl[7064], bl[7065], bl[7066], bl[7067], bl[7068], bl[7069], bl[7070], bl[7071], bl[7072], bl[7073], bl[7074], bl[7075], bl[7076], bl[7077], bl[7078], bl[7079], bl[7080], bl[7081], bl[7082], bl[7083], bl[7084], bl[7085], bl[7086], bl[7087], bl[7088], bl[7089], bl[7090], bl[7091], bl[7092], bl[7093], bl[7094], bl[7095], bl[7096], bl[7097], bl[7098], bl[7099], bl[7100], bl[7101], bl[7102], bl[7103], bl[7104], bl[7105], bl[7106], bl[7107], bl[7108], bl[7109], bl[7110], bl[7111], bl[7112], bl[7113], bl[7114], bl[7115], bl[7116], bl[7117], bl[7118], bl[7119], bl[7120], bl[7121], bl[7122], bl[7123], bl[7124], bl[7125], bl[7126], bl[7127], bl[7128], bl[7129], bl[7130], bl[7131], bl[7132], bl[7133], bl[7134], bl[7135], bl[7136], bl[7137], bl[7138], bl[7139], bl[7140], bl[7141], bl[7142], bl[7143], bl[7144], bl[7145], bl[7146], bl[7147], bl[7148], bl[7149], bl[7150], bl[7151], bl[7152], bl[7153], bl[7154], bl[7155], bl[7156], bl[7157], bl[7158], bl[7159], bl[7160], bl[7161], bl[7162], bl[7163], bl[7164], bl[7165], bl[7166], bl[7167], bl[7168], bl[7169], bl[7170], bl[7171], bl[7172], bl[7173], bl[7174], bl[7175], bl[7176], bl[7177], bl[7178], bl[7179], bl[7180], bl[7181], bl[7182], bl[7183], bl[7184], bl[7185], bl[7186], bl[7187], bl[7188], bl[7189], bl[7190], bl[7191], bl[7192], bl[7193], bl[7194], bl[7195], bl[7196], bl[7197], bl[7198], bl[7199], bl[7200], bl[7201], bl[7202], bl[7203], bl[7204], bl[7205], bl[7206], bl[7207], bl[7208], bl[7209], bl[7210], bl[7211], bl[7212], bl[7213], bl[7214], bl[7215], bl[7216], bl[7217], bl[7218], bl[7219], bl[7220], bl[7221], bl[7222], bl[7223], bl[7224], bl[7225], bl[7226], bl[7227], bl[7228], bl[7229], bl[7230], bl[7231], bl[7232], bl[7233], bl[7234], bl[7235], bl[7236], bl[7237], bl[7238], bl[7239], bl[7240], bl[7241], bl[7242], bl[7243], bl[7244], bl[7245], bl[7246], bl[7247], bl[7248], bl[7249], bl[7250], bl[7251], bl[7252], bl[7253], bl[7254], bl[7255], bl[7256], bl[7257], bl[7258], bl[7259], bl[7260], bl[7261], bl[7262], bl[7263], bl[7264], bl[7265], bl[7266], bl[7267], bl[7268], bl[7269], bl[7270], bl[7271], bl[7272], bl[7273], bl[7274], bl[7275], bl[7276], bl[7277], bl[7278], bl[7279], bl[7280], bl[7281], bl[7282], bl[7283], bl[7284], bl[7285], bl[7286], bl[7287], bl[7288], bl[7289], bl[7290], bl[7291], bl[7292], bl[7293], bl[7294], bl[7295], bl[7296], bl[7297], bl[7298], bl[7299], bl[7300], bl[7301], bl[7302], bl[7303], bl[7304], bl[7305], bl[7306], bl[7307], bl[7308], bl[7309], bl[7310], bl[7311], bl[7312], bl[7313], bl[7314], bl[7315], bl[7316], bl[7317], bl[7318], bl[7319], bl[7320], bl[7321], bl[7322], bl[7323], bl[7324], bl[7325], bl[7326], bl[7327], bl[7328], bl[7329], bl[7330], bl[7331], bl[7332], bl[7333], bl[7334], bl[7335], bl[7336], bl[7337], bl[7338], bl[7339], bl[7340], bl[7341], bl[7342], bl[7343], bl[7344], bl[7345], bl[7346], bl[7347], bl[7348], bl[7349], bl[7350], bl[7351], bl[7352], bl[7353], bl[7354], bl[7355], bl[7356], bl[7357], bl[7358], bl[7359], bl[7360], bl[7361], bl[7362], bl[7363], bl[7364], bl[7365], bl[7366], bl[7367], bl[7368], bl[7369], bl[7370], bl[7371], bl[7372], bl[7373], bl[7374], bl[7375], bl[7376], bl[7377], bl[7378], bl[7379], bl[7380], bl[7381], bl[7382], bl[7383], bl[7384], bl[7385], bl[7386], bl[7387], bl[7388], bl[7389], bl[7390], bl[7391], bl[7392], bl[7393], bl[7394], bl[7395], bl[7396], bl[7397], bl[7398], bl[7399], bl[7400], bl[7401], bl[7402], bl[7403], bl[7404], bl[7405], bl[7406], bl[7407], bl[7408], bl[7409], bl[7410], bl[7411], bl[7412], bl[7413], bl[7414], bl[7415], bl[7416], bl[7417], bl[7418], bl[7419], bl[7420], bl[7421], bl[7422], bl[7423], bl[7424], bl[7425], bl[7426], bl[7427], bl[7428], bl[7429], bl[7430], bl[7431], bl[7432], bl[7433], bl[7434], bl[7435], bl[7436], bl[7437], bl[7438], bl[7439], bl[7440], bl[7441], bl[7442], bl[7443], bl[7444], bl[7445], bl[7446], bl[7447], bl[7448], bl[7449], bl[7450], bl[7451], bl[7452], bl[7453], bl[7454], bl[7455], bl[7456], bl[7457], bl[7458], bl[7459], bl[7460], bl[7461], bl[7462], bl[7463], bl[7464], bl[7465], bl[7466], bl[7467], bl[7468], bl[7469], bl[7470], bl[7471], bl[7472], bl[7473], bl[7474], bl[7475], bl[7476], bl[7477], bl[7478], bl[7479], bl[7480], bl[7481], bl[7482], bl[7483], bl[7484], bl[7485], bl[7486], bl[7487], bl[7488], bl[7489], bl[7490], bl[7491], bl[7492], bl[7493], bl[7494], bl[7495], bl[7496], bl[7497], bl[7498], bl[7499], bl[7500], bl[7501], bl[7502], bl[7503], bl[7504], bl[7505], bl[7506], bl[7507], bl[7508], bl[7509], bl[7510], bl[7511], bl[7512], bl[7513], bl[7514], bl[7515], bl[7516], bl[7517], bl[7518], bl[7519], bl[7520], bl[7521], bl[7522], bl[7523], bl[7524], bl[7525], bl[7526], bl[7527], bl[7528], bl[7529], bl[7530], bl[7531], bl[7532], bl[7533], bl[7534], bl[7535], bl[7536], bl[7537], bl[7538], bl[7539], bl[7540], bl[7541], bl[7542], bl[7543], bl[7544], bl[7545], bl[7546], bl[7547], bl[7548], bl[7549], bl[7550], bl[7551], bl[7552], bl[7553], bl[7554], bl[7555], bl[7556], bl[7557], bl[7558], bl[7559], bl[7560], bl[7561], bl[7562], bl[7563], bl[7564], bl[7565], bl[7566], bl[7567], bl[7568], bl[7569], bl[7570], bl[7571], bl[7572], bl[7573], bl[7574], bl[7575], bl[7576], bl[7577], bl[7578], bl[7579], bl[7580], bl[7581], bl[7582], bl[7583], bl[7584], bl[7585], bl[7586], bl[7587], bl[7588], bl[7589], bl[7590], bl[7591], bl[7592], bl[7593], bl[7594], bl[7595], bl[7596], bl[7597], bl[7598], bl[7599], bl[7600], bl[7601], bl[7602], bl[7603], bl[7604], bl[7605], bl[7606], bl[7607], bl[7608], bl[7609], bl[7610], bl[7611], bl[7612], bl[7613], bl[7614], bl[7615], bl[7616], bl[7617], bl[7618], bl[7619], bl[7620], bl[7621], bl[7622], bl[7623], bl[7624], bl[7625], bl[7626], bl[7627], bl[7628], bl[7629], bl[7630], bl[7631], bl[7632], bl[7633], bl[7634], bl[7635], bl[7636], bl[7637], bl[7638], bl[7639], bl[7640], bl[7641], bl[7642], bl[7643], bl[7644], bl[7645], bl[7646], bl[7647], bl[7648], bl[7649], bl[7650], bl[7651], bl[7652], bl[7653], bl[7654], bl[7655], bl[7656], bl[7657], bl[7658], bl[7659], bl[7660], bl[7661], bl[7662], bl[7663], bl[15304], bl[15305], bl[15306], bl[15307], bl[15308], bl[15309], bl[15310], bl[15311], bl[15312], bl[15313], bl[15314], bl[15315], bl[15316], bl[15317], bl[15318], bl[15319], bl[15320], bl[15321], bl[15322], bl[15323], bl[15324], bl[15325], bl[15326], bl[15327], bl[15328], bl[15329], bl[15330], bl[15331], bl[15332], bl[15333], bl[15334], bl[15335], bl[15336], bl[15337], bl[15338], bl[15339], bl[15340], bl[15341], bl[15342], bl[15343], bl[15344], bl[15345], bl[15346], bl[15347], bl[15348], bl[15349], bl[15350], bl[15351], bl[15352], bl[15353], bl[15354], bl[15355], bl[15356], bl[15357], bl[15358], bl[15359], bl[15360], bl[15361], bl[15362], bl[15363], bl[15364], bl[15365], bl[15366], bl[15367], bl[15368], bl[15369], bl[15370], bl[15371], bl[15372], bl[15373], bl[15374], bl[15375], bl[15376], bl[15377], bl[15378], bl[15379], bl[15380], bl[15381], bl[15382], bl[15383], bl[40], bl[41], bl[42], bl[43], bl[44], bl[45], bl[46], bl[47], bl[6572], bl[6573], bl[6574], bl[6575], bl[6576], bl[6577], bl[6578], bl[6579], bl[6580], bl[6581], bl[6582], bl[6583], bl[6584], bl[6585], bl[6586], bl[6587], bl[6588], bl[6589], bl[6590], bl[6591], bl[6592], bl[6593], bl[6594], bl[6595], bl[6596], bl[6597], bl[6598], bl[6599], bl[6600], bl[6601], bl[6602], bl[6603], bl[6604], bl[6605], bl[6606], bl[6607], bl[6608], bl[6609], bl[6610], bl[6611], bl[6612], bl[6613], bl[6614], bl[6615], bl[6616], bl[6617], bl[6618], bl[6619], bl[6620], bl[6621], bl[6622], bl[6623], bl[6624], bl[6625], bl[6626], bl[6627], bl[6628], bl[6629], bl[6630], bl[6631], bl[6632], bl[6633], bl[6634], bl[6635], bl[6636], bl[6637], bl[6638], bl[6639], bl[6640], bl[6641], bl[6642], bl[6643], bl[15224], bl[15225], bl[15226], bl[15227], bl[15228], bl[15229], bl[15230], bl[15231], bl[15232], bl[15233], bl[15234], bl[15235], bl[15236], bl[15237], bl[15238], bl[15239], bl[15240], bl[15241], bl[15242], bl[15243], bl[15244], bl[15245], bl[15246], bl[15247], bl[15248], bl[15249], bl[15250], bl[15251], bl[15252], bl[15253], bl[15254], bl[15255], bl[15256], bl[15257], bl[15258], bl[15259], bl[15260], bl[15261], bl[15262], bl[15263], bl[15264], bl[15265], bl[15266], bl[15267], bl[15268], bl[15269], bl[15270], bl[15271], bl[15272], bl[15273], bl[15274], bl[15275], bl[15276], bl[15277], bl[15278], bl[15279], bl[15280], bl[15281], bl[15282], bl[15283], bl[15284], bl[15285], bl[15286], bl[15287], bl[15288], bl[15289], bl[15290], bl[15291], bl[15292], bl[15293], bl[15294], bl[15295], bl[15296], bl[15297], bl[15298], bl[15299], bl[15300], bl[15301], bl[15302], bl[15303]}),
        .wl({wl[6644], wl[6645], wl[6646], wl[6647], wl[6648], wl[6649], wl[6650], wl[6651], wl[6652], wl[6653], wl[6654], wl[6655], wl[6656], wl[6657], wl[6658], wl[6659], wl[6660], wl[6661], wl[6662], wl[6663], wl[6664], wl[6665], wl[6666], wl[6667], wl[6668], wl[6669], wl[6670], wl[6671], wl[6672], wl[6673], wl[6674], wl[6675], wl[6676], wl[6677], wl[6678], wl[6679], wl[6680], wl[6681], wl[6682], wl[6683], wl[6684], wl[6685], wl[6686], wl[6687], wl[6688], wl[6689], wl[6690], wl[6691], wl[6692], wl[6693], wl[6694], wl[6695], wl[6696], wl[6697], wl[6698], wl[6699], wl[6700], wl[6701], wl[6702], wl[6703], wl[6704], wl[6705], wl[6706], wl[6707], wl[6708], wl[6709], wl[6710], wl[6711], wl[6712], wl[6713], wl[6714], wl[6715], wl[6716], wl[6717], wl[6718], wl[6719], wl[6720], wl[6721], wl[6722], wl[6723], wl[6724], wl[6725], wl[6726], wl[6727], wl[6728], wl[6729], wl[6730], wl[6731], wl[6732], wl[6733], wl[6734], wl[6735], wl[6736], wl[6737], wl[6738], wl[6739], wl[6740], wl[6741], wl[6742], wl[6743], wl[6744], wl[6745], wl[6746], wl[6747], wl[6748], wl[6749], wl[6750], wl[6751], wl[6752], wl[6753], wl[6754], wl[6755], wl[6756], wl[6757], wl[6758], wl[6759], wl[6760], wl[6761], wl[6762], wl[6763], wl[6764], wl[6765], wl[6766], wl[6767], wl[6768], wl[6769], wl[6770], wl[6771], wl[6772], wl[6773], wl[6774], wl[6775], wl[6776], wl[6777], wl[6778], wl[6779], wl[6780], wl[6781], wl[6782], wl[6783], wl[6784], wl[6785], wl[6786], wl[6787], wl[6788], wl[6789], wl[6790], wl[6791], wl[6792], wl[6793], wl[6794], wl[6795], wl[6796], wl[6797], wl[6798], wl[6799], wl[6800], wl[6801], wl[6802], wl[6803], wl[6804], wl[6805], wl[6806], wl[6807], wl[6808], wl[6809], wl[6810], wl[6811], wl[6812], wl[6813], wl[6814], wl[6815], wl[6816], wl[6817], wl[6818], wl[6819], wl[6820], wl[6821], wl[6822], wl[6823], wl[6824], wl[6825], wl[6826], wl[6827], wl[6828], wl[6829], wl[6830], wl[6831], wl[6832], wl[6833], wl[6834], wl[6835], wl[6836], wl[6837], wl[6838], wl[6839], wl[6840], wl[6841], wl[6842], wl[6843], wl[6844], wl[6845], wl[6846], wl[6847], wl[6848], wl[6849], wl[6850], wl[6851], wl[6852], wl[6853], wl[6854], wl[6855], wl[6856], wl[6857], wl[6858], wl[6859], wl[6860], wl[6861], wl[6862], wl[6863], wl[6864], wl[6865], wl[6866], wl[6867], wl[6868], wl[6869], wl[6870], wl[6871], wl[6872], wl[6873], wl[6874], wl[6875], wl[6876], wl[6877], wl[6878], wl[6879], wl[6880], wl[6881], wl[6882], wl[6883], wl[6884], wl[6885], wl[6886], wl[6887], wl[6888], wl[6889], wl[6890], wl[6891], wl[6892], wl[6893], wl[6894], wl[6895], wl[6896], wl[6897], wl[6898], wl[6899], wl[6900], wl[6901], wl[6902], wl[6903], wl[6904], wl[6905], wl[6906], wl[6907], wl[6908], wl[6909], wl[6910], wl[6911], wl[6912], wl[6913], wl[6914], wl[6915], wl[6916], wl[6917], wl[6918], wl[6919], wl[6920], wl[6921], wl[6922], wl[6923], wl[6924], wl[6925], wl[6926], wl[6927], wl[6928], wl[6929], wl[6930], wl[6931], wl[6932], wl[6933], wl[6934], wl[6935], wl[6936], wl[6937], wl[6938], wl[6939], wl[6940], wl[6941], wl[6942], wl[6943], wl[6944], wl[6945], wl[6946], wl[6947], wl[6948], wl[6949], wl[6950], wl[6951], wl[6952], wl[6953], wl[6954], wl[6955], wl[6956], wl[6957], wl[6958], wl[6959], wl[6960], wl[6961], wl[6962], wl[6963], wl[6964], wl[6965], wl[6966], wl[6967], wl[6968], wl[6969], wl[6970], wl[6971], wl[6972], wl[6973], wl[6974], wl[6975], wl[6976], wl[6977], wl[6978], wl[6979], wl[6980], wl[6981], wl[6982], wl[6983], wl[6984], wl[6985], wl[6986], wl[6987], wl[6988], wl[6989], wl[6990], wl[6991], wl[6992], wl[6993], wl[6994], wl[6995], wl[6996], wl[6997], wl[6998], wl[6999], wl[7000], wl[7001], wl[7002], wl[7003], wl[7004], wl[7005], wl[7006], wl[7007], wl[7008], wl[7009], wl[7010], wl[7011], wl[7012], wl[7013], wl[7014], wl[7015], wl[7016], wl[7017], wl[7018], wl[7019], wl[7020], wl[7021], wl[7022], wl[7023], wl[7024], wl[7025], wl[7026], wl[7027], wl[7028], wl[7029], wl[7030], wl[7031], wl[7032], wl[7033], wl[7034], wl[7035], wl[7036], wl[7037], wl[7038], wl[7039], wl[7040], wl[7041], wl[7042], wl[7043], wl[7044], wl[7045], wl[7046], wl[7047], wl[7048], wl[7049], wl[7050], wl[7051], wl[7052], wl[7053], wl[7054], wl[7055], wl[7056], wl[7057], wl[7058], wl[7059], wl[7060], wl[7061], wl[7062], wl[7063], wl[7064], wl[7065], wl[7066], wl[7067], wl[7068], wl[7069], wl[7070], wl[7071], wl[7072], wl[7073], wl[7074], wl[7075], wl[7076], wl[7077], wl[7078], wl[7079], wl[7080], wl[7081], wl[7082], wl[7083], wl[7084], wl[7085], wl[7086], wl[7087], wl[7088], wl[7089], wl[7090], wl[7091], wl[7092], wl[7093], wl[7094], wl[7095], wl[7096], wl[7097], wl[7098], wl[7099], wl[7100], wl[7101], wl[7102], wl[7103], wl[7104], wl[7105], wl[7106], wl[7107], wl[7108], wl[7109], wl[7110], wl[7111], wl[7112], wl[7113], wl[7114], wl[7115], wl[7116], wl[7117], wl[7118], wl[7119], wl[7120], wl[7121], wl[7122], wl[7123], wl[7124], wl[7125], wl[7126], wl[7127], wl[7128], wl[7129], wl[7130], wl[7131], wl[7132], wl[7133], wl[7134], wl[7135], wl[7136], wl[7137], wl[7138], wl[7139], wl[7140], wl[7141], wl[7142], wl[7143], wl[7144], wl[7145], wl[7146], wl[7147], wl[7148], wl[7149], wl[7150], wl[7151], wl[7152], wl[7153], wl[7154], wl[7155], wl[7156], wl[7157], wl[7158], wl[7159], wl[7160], wl[7161], wl[7162], wl[7163], wl[7164], wl[7165], wl[7166], wl[7167], wl[7168], wl[7169], wl[7170], wl[7171], wl[7172], wl[7173], wl[7174], wl[7175], wl[7176], wl[7177], wl[7178], wl[7179], wl[7180], wl[7181], wl[7182], wl[7183], wl[7184], wl[7185], wl[7186], wl[7187], wl[7188], wl[7189], wl[7190], wl[7191], wl[7192], wl[7193], wl[7194], wl[7195], wl[7196], wl[7197], wl[7198], wl[7199], wl[7200], wl[7201], wl[7202], wl[7203], wl[7204], wl[7205], wl[7206], wl[7207], wl[7208], wl[7209], wl[7210], wl[7211], wl[7212], wl[7213], wl[7214], wl[7215], wl[7216], wl[7217], wl[7218], wl[7219], wl[7220], wl[7221], wl[7222], wl[7223], wl[7224], wl[7225], wl[7226], wl[7227], wl[7228], wl[7229], wl[7230], wl[7231], wl[7232], wl[7233], wl[7234], wl[7235], wl[7236], wl[7237], wl[7238], wl[7239], wl[7240], wl[7241], wl[7242], wl[7243], wl[7244], wl[7245], wl[7246], wl[7247], wl[7248], wl[7249], wl[7250], wl[7251], wl[7252], wl[7253], wl[7254], wl[7255], wl[7256], wl[7257], wl[7258], wl[7259], wl[7260], wl[7261], wl[7262], wl[7263], wl[7264], wl[7265], wl[7266], wl[7267], wl[7268], wl[7269], wl[7270], wl[7271], wl[7272], wl[7273], wl[7274], wl[7275], wl[7276], wl[7277], wl[7278], wl[7279], wl[7280], wl[7281], wl[7282], wl[7283], wl[7284], wl[7285], wl[7286], wl[7287], wl[7288], wl[7289], wl[7290], wl[7291], wl[7292], wl[7293], wl[7294], wl[7295], wl[7296], wl[7297], wl[7298], wl[7299], wl[7300], wl[7301], wl[7302], wl[7303], wl[7304], wl[7305], wl[7306], wl[7307], wl[7308], wl[7309], wl[7310], wl[7311], wl[7312], wl[7313], wl[7314], wl[7315], wl[7316], wl[7317], wl[7318], wl[7319], wl[7320], wl[7321], wl[7322], wl[7323], wl[7324], wl[7325], wl[7326], wl[7327], wl[7328], wl[7329], wl[7330], wl[7331], wl[7332], wl[7333], wl[7334], wl[7335], wl[7336], wl[7337], wl[7338], wl[7339], wl[7340], wl[7341], wl[7342], wl[7343], wl[7344], wl[7345], wl[7346], wl[7347], wl[7348], wl[7349], wl[7350], wl[7351], wl[7352], wl[7353], wl[7354], wl[7355], wl[7356], wl[7357], wl[7358], wl[7359], wl[7360], wl[7361], wl[7362], wl[7363], wl[7364], wl[7365], wl[7366], wl[7367], wl[7368], wl[7369], wl[7370], wl[7371], wl[7372], wl[7373], wl[7374], wl[7375], wl[7376], wl[7377], wl[7378], wl[7379], wl[7380], wl[7381], wl[7382], wl[7383], wl[7384], wl[7385], wl[7386], wl[7387], wl[7388], wl[7389], wl[7390], wl[7391], wl[7392], wl[7393], wl[7394], wl[7395], wl[7396], wl[7397], wl[7398], wl[7399], wl[7400], wl[7401], wl[7402], wl[7403], wl[7404], wl[7405], wl[7406], wl[7407], wl[7408], wl[7409], wl[7410], wl[7411], wl[7412], wl[7413], wl[7414], wl[7415], wl[7416], wl[7417], wl[7418], wl[7419], wl[7420], wl[7421], wl[7422], wl[7423], wl[7424], wl[7425], wl[7426], wl[7427], wl[7428], wl[7429], wl[7430], wl[7431], wl[7432], wl[7433], wl[7434], wl[7435], wl[7436], wl[7437], wl[7438], wl[7439], wl[7440], wl[7441], wl[7442], wl[7443], wl[7444], wl[7445], wl[7446], wl[7447], wl[7448], wl[7449], wl[7450], wl[7451], wl[7452], wl[7453], wl[7454], wl[7455], wl[7456], wl[7457], wl[7458], wl[7459], wl[7460], wl[7461], wl[7462], wl[7463], wl[7464], wl[7465], wl[7466], wl[7467], wl[7468], wl[7469], wl[7470], wl[7471], wl[7472], wl[7473], wl[7474], wl[7475], wl[7476], wl[7477], wl[7478], wl[7479], wl[7480], wl[7481], wl[7482], wl[7483], wl[7484], wl[7485], wl[7486], wl[7487], wl[7488], wl[7489], wl[7490], wl[7491], wl[7492], wl[7493], wl[7494], wl[7495], wl[7496], wl[7497], wl[7498], wl[7499], wl[7500], wl[7501], wl[7502], wl[7503], wl[7504], wl[7505], wl[7506], wl[7507], wl[7508], wl[7509], wl[7510], wl[7511], wl[7512], wl[7513], wl[7514], wl[7515], wl[7516], wl[7517], wl[7518], wl[7519], wl[7520], wl[7521], wl[7522], wl[7523], wl[7524], wl[7525], wl[7526], wl[7527], wl[7528], wl[7529], wl[7530], wl[7531], wl[7532], wl[7533], wl[7534], wl[7535], wl[7536], wl[7537], wl[7538], wl[7539], wl[7540], wl[7541], wl[7542], wl[7543], wl[7544], wl[7545], wl[7546], wl[7547], wl[7548], wl[7549], wl[7550], wl[7551], wl[7552], wl[7553], wl[7554], wl[7555], wl[7556], wl[7557], wl[7558], wl[7559], wl[7560], wl[7561], wl[7562], wl[7563], wl[7564], wl[7565], wl[7566], wl[7567], wl[7568], wl[7569], wl[7570], wl[7571], wl[7572], wl[7573], wl[7574], wl[7575], wl[7576], wl[7577], wl[7578], wl[7579], wl[7580], wl[7581], wl[7582], wl[7583], wl[7584], wl[7585], wl[7586], wl[7587], wl[7588], wl[7589], wl[7590], wl[7591], wl[7592], wl[7593], wl[7594], wl[7595], wl[7596], wl[7597], wl[7598], wl[7599], wl[7600], wl[7601], wl[7602], wl[7603], wl[7604], wl[7605], wl[7606], wl[7607], wl[7608], wl[7609], wl[7610], wl[7611], wl[7612], wl[7613], wl[7614], wl[7615], wl[7616], wl[7617], wl[7618], wl[7619], wl[7620], wl[7621], wl[7622], wl[7623], wl[7624], wl[7625], wl[7626], wl[7627], wl[7628], wl[7629], wl[7630], wl[7631], wl[7632], wl[7633], wl[7634], wl[7635], wl[7636], wl[7637], wl[7638], wl[7639], wl[7640], wl[7641], wl[7642], wl[7643], wl[7644], wl[7645], wl[7646], wl[7647], wl[7648], wl[7649], wl[7650], wl[7651], wl[7652], wl[7653], wl[7654], wl[7655], wl[7656], wl[7657], wl[7658], wl[7659], wl[7660], wl[7661], wl[7662], wl[7663], wl[15304], wl[15305], wl[15306], wl[15307], wl[15308], wl[15309], wl[15310], wl[15311], wl[15312], wl[15313], wl[15314], wl[15315], wl[15316], wl[15317], wl[15318], wl[15319], wl[15320], wl[15321], wl[15322], wl[15323], wl[15324], wl[15325], wl[15326], wl[15327], wl[15328], wl[15329], wl[15330], wl[15331], wl[15332], wl[15333], wl[15334], wl[15335], wl[15336], wl[15337], wl[15338], wl[15339], wl[15340], wl[15341], wl[15342], wl[15343], wl[15344], wl[15345], wl[15346], wl[15347], wl[15348], wl[15349], wl[15350], wl[15351], wl[15352], wl[15353], wl[15354], wl[15355], wl[15356], wl[15357], wl[15358], wl[15359], wl[15360], wl[15361], wl[15362], wl[15363], wl[15364], wl[15365], wl[15366], wl[15367], wl[15368], wl[15369], wl[15370], wl[15371], wl[15372], wl[15373], wl[15374], wl[15375], wl[15376], wl[15377], wl[15378], wl[15379], wl[15380], wl[15381], wl[15382], wl[15383], wl[40], wl[41], wl[42], wl[43], wl[44], wl[45], wl[46], wl[47], wl[6572], wl[6573], wl[6574], wl[6575], wl[6576], wl[6577], wl[6578], wl[6579], wl[6580], wl[6581], wl[6582], wl[6583], wl[6584], wl[6585], wl[6586], wl[6587], wl[6588], wl[6589], wl[6590], wl[6591], wl[6592], wl[6593], wl[6594], wl[6595], wl[6596], wl[6597], wl[6598], wl[6599], wl[6600], wl[6601], wl[6602], wl[6603], wl[6604], wl[6605], wl[6606], wl[6607], wl[6608], wl[6609], wl[6610], wl[6611], wl[6612], wl[6613], wl[6614], wl[6615], wl[6616], wl[6617], wl[6618], wl[6619], wl[6620], wl[6621], wl[6622], wl[6623], wl[6624], wl[6625], wl[6626], wl[6627], wl[6628], wl[6629], wl[6630], wl[6631], wl[6632], wl[6633], wl[6634], wl[6635], wl[6636], wl[6637], wl[6638], wl[6639], wl[6640], wl[6641], wl[6642], wl[6643], wl[15224], wl[15225], wl[15226], wl[15227], wl[15228], wl[15229], wl[15230], wl[15231], wl[15232], wl[15233], wl[15234], wl[15235], wl[15236], wl[15237], wl[15238], wl[15239], wl[15240], wl[15241], wl[15242], wl[15243], wl[15244], wl[15245], wl[15246], wl[15247], wl[15248], wl[15249], wl[15250], wl[15251], wl[15252], wl[15253], wl[15254], wl[15255], wl[15256], wl[15257], wl[15258], wl[15259], wl[15260], wl[15261], wl[15262], wl[15263], wl[15264], wl[15265], wl[15266], wl[15267], wl[15268], wl[15269], wl[15270], wl[15271], wl[15272], wl[15273], wl[15274], wl[15275], wl[15276], wl[15277], wl[15278], wl[15279], wl[15280], wl[15281], wl[15282], wl[15283], wl[15284], wl[15285], wl[15286], wl[15287], wl[15288], wl[15289], wl[15290], wl[15291], wl[15292], wl[15293], wl[15294], wl[15295], wl[15296], wl[15297], wl[15298], wl[15299], wl[15300], wl[15301], wl[15302], wl[15303]})
    );
    right_tile tile_5__4_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_3__3__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_3__3__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_3__3__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_4__2__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_4__2__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_4__2__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_3__2__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_3__2__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_3__2__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_3__2__grid_top_r_in[1]),
        .grid_left_in(grid_clb_4__3__grid_left_in),
        .grid_bottom_in(grid_clb_4__3__grid_bottom_in),
        .chanx_left_in(sb_1__1__8_chanx_right_out),
        .chanx_left_out(cbx_1__1__11_chanx_left_out),
        .grid_top_out(grid_clb_4__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[40:47]),
        .io_left_in(grid_io_right_5__3__io_left_in),
        .chany_bottom_in(sb_4__1__1_chany_top_out),
        .chany_bottom_out(cby_4__1__2_chany_bottom_out),
        .chany_top_in_0(cby_4__1__3_chany_bottom_out),
        .chany_top_out_0(sb_4__1__2_chany_top_out),
        .grid_top_r_inpad(grid_io_right_5__4__io_left_in),
        .grid_top_l_in(sb_4__3__grid_top_l_in),
        .grid_bottom_l_in(sb_4__2__grid_top_l_in),
        .grid_left_t_in(sb_3__3__grid_right_t_in),
        .grid_left_b_in(sb_3__3__grid_right_b_in),
        .bl({bl[15456], bl[15457], bl[15458], bl[15459], bl[15460], bl[15461], bl[15462], bl[15463], bl[15464], bl[15465], bl[15466], bl[15467], bl[15468], bl[15469], bl[15470], bl[15471], bl[15472], bl[15473], bl[15474], bl[15475], bl[15476], bl[15477], bl[15478], bl[15479], bl[15480], bl[15481], bl[15482], bl[15483], bl[15484], bl[15485], bl[15486], bl[15487], bl[15488], bl[15489], bl[15490], bl[15491], bl[15492], bl[15493], bl[15494], bl[15495], bl[15496], bl[15497], bl[15498], bl[15499], bl[15500], bl[15501], bl[15502], bl[15503], bl[15504], bl[15505], bl[15506], bl[15507], bl[15508], bl[15509], bl[15510], bl[15511], bl[15512], bl[15513], bl[15514], bl[15515], bl[15516], bl[15517], bl[15518], bl[15519], bl[15520], bl[15521], bl[15522], bl[15523], bl[15524], bl[15525], bl[15526], bl[15527], bl[15528], bl[15529], bl[15530], bl[15531], bl[15532], bl[15533], bl[15534], bl[15535], bl[15536], bl[15537], bl[15538], bl[15539], bl[15540], bl[15541], bl[15542], bl[15543], bl[15544], bl[15545], bl[15546], bl[15547], bl[15548], bl[15549], bl[15550], bl[15551], bl[15552], bl[15553], bl[15554], bl[15555], bl[15556], bl[15557], bl[15558], bl[15559], bl[15560], bl[15561], bl[15562], bl[15563], bl[15564], bl[15565], bl[15566], bl[15567], bl[15568], bl[15569], bl[15570], bl[15571], bl[15572], bl[15573], bl[15574], bl[15575], bl[15576], bl[15577], bl[15578], bl[15579], bl[15580], bl[15581], bl[15582], bl[15583], bl[15584], bl[15585], bl[15586], bl[15587], bl[15588], bl[15589], bl[15590], bl[15591], bl[15592], bl[15593], bl[15594], bl[15595], bl[15596], bl[15597], bl[15598], bl[15599], bl[15600], bl[15601], bl[15602], bl[15603], bl[15604], bl[15605], bl[15606], bl[15607], bl[15608], bl[15609], bl[15610], bl[15611], bl[15612], bl[15613], bl[15614], bl[15615], bl[15616], bl[15617], bl[15618], bl[15619], bl[15620], bl[15621], bl[15622], bl[15623], bl[15624], bl[15625], bl[15626], bl[15627], bl[15628], bl[15629], bl[15630], bl[15631], bl[15632], bl[15633], bl[15634], bl[15635], bl[15636], bl[15637], bl[15638], bl[15639], bl[15640], bl[15641], bl[15642], bl[15643], bl[15644], bl[15645], bl[15646], bl[15647], bl[15648], bl[15649], bl[15650], bl[15651], bl[15652], bl[15653], bl[15654], bl[15655], bl[15656], bl[15657], bl[15658], bl[15659], bl[15660], bl[15661], bl[15662], bl[15663], bl[15664], bl[15665], bl[15666], bl[15667], bl[15668], bl[15669], bl[15670], bl[15671], bl[15672], bl[15673], bl[15674], bl[15675], bl[15676], bl[15677], bl[15678], bl[15679], bl[15680], bl[15681], bl[15682], bl[15683], bl[15684], bl[15685], bl[15686], bl[15687], bl[15688], bl[15689], bl[15690], bl[15691], bl[15692], bl[15693], bl[15694], bl[15695], bl[15696], bl[15697], bl[15698], bl[15699], bl[15700], bl[15701], bl[15702], bl[15703], bl[15704], bl[15705], bl[15706], bl[15707], bl[15708], bl[15709], bl[15710], bl[15711], bl[15712], bl[15713], bl[15714], bl[15715], bl[15716], bl[15717], bl[15718], bl[15719], bl[15720], bl[15721], bl[15722], bl[15723], bl[15724], bl[15725], bl[15726], bl[15727], bl[15728], bl[15729], bl[15730], bl[15731], bl[15732], bl[15733], bl[15734], bl[15735], bl[15736], bl[15737], bl[15738], bl[15739], bl[15740], bl[15741], bl[15742], bl[15743], bl[15744], bl[15745], bl[15746], bl[15747], bl[15748], bl[15749], bl[15750], bl[15751], bl[15752], bl[15753], bl[15754], bl[15755], bl[15756], bl[15757], bl[15758], bl[15759], bl[15760], bl[15761], bl[15762], bl[15763], bl[15764], bl[15765], bl[15766], bl[15767], bl[15768], bl[15769], bl[15770], bl[15771], bl[15772], bl[15773], bl[15774], bl[15775], bl[15776], bl[15777], bl[15778], bl[15779], bl[15780], bl[15781], bl[15782], bl[15783], bl[15784], bl[15785], bl[15786], bl[15787], bl[15788], bl[15789], bl[15790], bl[15791], bl[15792], bl[15793], bl[15794], bl[15795], bl[15796], bl[15797], bl[15798], bl[15799], bl[15800], bl[15801], bl[15802], bl[15803], bl[15804], bl[15805], bl[15806], bl[15807], bl[15808], bl[15809], bl[15810], bl[15811], bl[15812], bl[15813], bl[15814], bl[15815], bl[15816], bl[15817], bl[15818], bl[15819], bl[15820], bl[15821], bl[15822], bl[15823], bl[15824], bl[15825], bl[15826], bl[15827], bl[15828], bl[15829], bl[15830], bl[15831], bl[15832], bl[15833], bl[15834], bl[15835], bl[15836], bl[15837], bl[15838], bl[15839], bl[15840], bl[15841], bl[15842], bl[15843], bl[15844], bl[15845], bl[15846], bl[15847], bl[15848], bl[15849], bl[15850], bl[15851], bl[15852], bl[15853], bl[15854], bl[15855], bl[15856], bl[15857], bl[15858], bl[15859], bl[15860], bl[15861], bl[15862], bl[15863], bl[15864], bl[15865], bl[15866], bl[15867], bl[15868], bl[15869], bl[15870], bl[15871], bl[15872], bl[15873], bl[15874], bl[15875], bl[15876], bl[15877], bl[15878], bl[15879], bl[15880], bl[15881], bl[15882], bl[15883], bl[15884], bl[15885], bl[15886], bl[15887], bl[15888], bl[15889], bl[15890], bl[15891], bl[15892], bl[15893], bl[15894], bl[15895], bl[15896], bl[15897], bl[15898], bl[15899], bl[15900], bl[15901], bl[15902], bl[15903], bl[15904], bl[15905], bl[15906], bl[15907], bl[15908], bl[15909], bl[15910], bl[15911], bl[15912], bl[15913], bl[15914], bl[15915], bl[15916], bl[15917], bl[15918], bl[15919], bl[15920], bl[15921], bl[15922], bl[15923], bl[15924], bl[15925], bl[15926], bl[15927], bl[15928], bl[15929], bl[15930], bl[15931], bl[15932], bl[15933], bl[15934], bl[15935], bl[15936], bl[15937], bl[15938], bl[15939], bl[15940], bl[15941], bl[15942], bl[15943], bl[15944], bl[15945], bl[15946], bl[15947], bl[15948], bl[15949], bl[15950], bl[15951], bl[15952], bl[15953], bl[15954], bl[15955], bl[15956], bl[15957], bl[15958], bl[15959], bl[15960], bl[15961], bl[15962], bl[15963], bl[15964], bl[15965], bl[15966], bl[15967], bl[15968], bl[15969], bl[15970], bl[15971], bl[15972], bl[15973], bl[15974], bl[15975], bl[15976], bl[15977], bl[15978], bl[15979], bl[15980], bl[15981], bl[15982], bl[15983], bl[15984], bl[15985], bl[15986], bl[15987], bl[15988], bl[15989], bl[15990], bl[15991], bl[15992], bl[15993], bl[15994], bl[15995], bl[15996], bl[15997], bl[15998], bl[15999], bl[16000], bl[16001], bl[16002], bl[16003], bl[16004], bl[16005], bl[16006], bl[16007], bl[16008], bl[16009], bl[16010], bl[16011], bl[16012], bl[16013], bl[16014], bl[16015], bl[16016], bl[16017], bl[16018], bl[16019], bl[16020], bl[16021], bl[16022], bl[16023], bl[16024], bl[16025], bl[16026], bl[16027], bl[16028], bl[16029], bl[16030], bl[16031], bl[16032], bl[16033], bl[16034], bl[16035], bl[16036], bl[16037], bl[16038], bl[16039], bl[16040], bl[16041], bl[16042], bl[16043], bl[16044], bl[16045], bl[16046], bl[16047], bl[16048], bl[16049], bl[16050], bl[16051], bl[16052], bl[16053], bl[16054], bl[16055], bl[16056], bl[16057], bl[16058], bl[16059], bl[16060], bl[16061], bl[16062], bl[16063], bl[16064], bl[16065], bl[16066], bl[16067], bl[16068], bl[16069], bl[16070], bl[16071], bl[16072], bl[16073], bl[16074], bl[16075], bl[16076], bl[16077], bl[16078], bl[16079], bl[16080], bl[16081], bl[16082], bl[16083], bl[16084], bl[16085], bl[16086], bl[16087], bl[16088], bl[16089], bl[16090], bl[16091], bl[16092], bl[16093], bl[16094], bl[16095], bl[16096], bl[16097], bl[16098], bl[16099], bl[16100], bl[16101], bl[16102], bl[16103], bl[16104], bl[16105], bl[16106], bl[16107], bl[16108], bl[16109], bl[16110], bl[16111], bl[16112], bl[16113], bl[16114], bl[16115], bl[16116], bl[16117], bl[16118], bl[16119], bl[16120], bl[16121], bl[16122], bl[16123], bl[16124], bl[16125], bl[16126], bl[16127], bl[16128], bl[16129], bl[16130], bl[16131], bl[16132], bl[16133], bl[16134], bl[16135], bl[16136], bl[16137], bl[16138], bl[16139], bl[16140], bl[16141], bl[16142], bl[16143], bl[16144], bl[16145], bl[16146], bl[16147], bl[16148], bl[16149], bl[16150], bl[16151], bl[16152], bl[16153], bl[16154], bl[16155], bl[16156], bl[16157], bl[16158], bl[16159], bl[16160], bl[16161], bl[16162], bl[16163], bl[16164], bl[16165], bl[16166], bl[16167], bl[16168], bl[16169], bl[16170], bl[16171], bl[16172], bl[16173], bl[16174], bl[16175], bl[16176], bl[16177], bl[16178], bl[16179], bl[16180], bl[16181], bl[16182], bl[16183], bl[16184], bl[16185], bl[16186], bl[16187], bl[16188], bl[16189], bl[16190], bl[16191], bl[16192], bl[16193], bl[16194], bl[16195], bl[16196], bl[16197], bl[16198], bl[16199], bl[16200], bl[16201], bl[16202], bl[16203], bl[16204], bl[16205], bl[16206], bl[16207], bl[16208], bl[16209], bl[16210], bl[16211], bl[16212], bl[16213], bl[16214], bl[16215], bl[16216], bl[16217], bl[16218], bl[16219], bl[16220], bl[16221], bl[16222], bl[16223], bl[16224], bl[16225], bl[16226], bl[16227], bl[16228], bl[16229], bl[16230], bl[16231], bl[16232], bl[16233], bl[16234], bl[16235], bl[16236], bl[16237], bl[16238], bl[16239], bl[16240], bl[16241], bl[16242], bl[16243], bl[16244], bl[16245], bl[16246], bl[16247], bl[16248], bl[16249], bl[16250], bl[16251], bl[16252], bl[16253], bl[16254], bl[16255], bl[16256], bl[16257], bl[16258], bl[16259], bl[16260], bl[16261], bl[16262], bl[16263], bl[16264], bl[16265], bl[16266], bl[16267], bl[16268], bl[16269], bl[16270], bl[16271], bl[16272], bl[16273], bl[16274], bl[16275], bl[16276], bl[16277], bl[16278], bl[16279], bl[16280], bl[16281], bl[16282], bl[16283], bl[16284], bl[16285], bl[16286], bl[16287], bl[16288], bl[16289], bl[16290], bl[16291], bl[16292], bl[16293], bl[16294], bl[16295], bl[16296], bl[16297], bl[16298], bl[16299], bl[16300], bl[16301], bl[16302], bl[16303], bl[16304], bl[16305], bl[16306], bl[16307], bl[16308], bl[16309], bl[16310], bl[16311], bl[16312], bl[16313], bl[16314], bl[16315], bl[16316], bl[16317], bl[16318], bl[16319], bl[16320], bl[16321], bl[16322], bl[16323], bl[16324], bl[16325], bl[16326], bl[16327], bl[16328], bl[16329], bl[16330], bl[16331], bl[16332], bl[16333], bl[16334], bl[16335], bl[16336], bl[16337], bl[16338], bl[16339], bl[16340], bl[16341], bl[16342], bl[16343], bl[16344], bl[16345], bl[16346], bl[16347], bl[16348], bl[16349], bl[16350], bl[16351], bl[16352], bl[16353], bl[16354], bl[16355], bl[16356], bl[16357], bl[16358], bl[16359], bl[16360], bl[16361], bl[16362], bl[16363], bl[16364], bl[16365], bl[16366], bl[16367], bl[16368], bl[16369], bl[16370], bl[16371], bl[16372], bl[16373], bl[16374], bl[16375], bl[16376], bl[16377], bl[16378], bl[16379], bl[16380], bl[16381], bl[16382], bl[16383], bl[16384], bl[16385], bl[16386], bl[16387], bl[16388], bl[16389], bl[16390], bl[16391], bl[16392], bl[16393], bl[16394], bl[16395], bl[16396], bl[16397], bl[16398], bl[16399], bl[16400], bl[16401], bl[16402], bl[16403], bl[16404], bl[16405], bl[16406], bl[16407], bl[16408], bl[16409], bl[16410], bl[16411], bl[16412], bl[16413], bl[16414], bl[16415], bl[16416], bl[16417], bl[16418], bl[16419], bl[16420], bl[16421], bl[16422], bl[16423], bl[16424], bl[16425], bl[16426], bl[16427], bl[16428], bl[16429], bl[16430], bl[16431], bl[16432], bl[16433], bl[16434], bl[16435], bl[16436], bl[16437], bl[16438], bl[16439], bl[16440], bl[16441], bl[16442], bl[16443], bl[16444], bl[16445], bl[16446], bl[16447], bl[16448], bl[16449], bl[16450], bl[16451], bl[16452], bl[16453], bl[16454], bl[16455], bl[16456], bl[16457], bl[16458], bl[16459], bl[16460], bl[16461], bl[16462], bl[16463], bl[16464], bl[16465], bl[16466], bl[16467], bl[16468], bl[16469], bl[16470], bl[16471], bl[16472], bl[16473], bl[16474], bl[16475], bl[16556], bl[16557], bl[16558], bl[16559], bl[16560], bl[16561], bl[16562], bl[16563], bl[16564], bl[16565], bl[16566], bl[16567], bl[16568], bl[16569], bl[16570], bl[16571], bl[16572], bl[16573], bl[16574], bl[16575], bl[16576], bl[16577], bl[16578], bl[16579], bl[16580], bl[16581], bl[16582], bl[16583], bl[16584], bl[16585], bl[16586], bl[16587], bl[16588], bl[16589], bl[16590], bl[16591], bl[16592], bl[16593], bl[16594], bl[16595], bl[16596], bl[16597], bl[16598], bl[16599], bl[16600], bl[16601], bl[16602], bl[16603], bl[16604], bl[16605], bl[16606], bl[16607], bl[16608], bl[16609], bl[16610], bl[16611], bl[16612], bl[16613], bl[16614], bl[16615], bl[16616], bl[16617], bl[16618], bl[16619], bl[16620], bl[16621], bl[16622], bl[16623], bl[16624], bl[16625], bl[16626], bl[16627], bl[16628], bl[16629], bl[16630], bl[16631], bl[16632], bl[16633], bl[16634], bl[16635], bl[48], bl[49], bl[50], bl[51], bl[52], bl[53], bl[54], bl[55], bl[15384], bl[15385], bl[15386], bl[15387], bl[15388], bl[15389], bl[15390], bl[15391], bl[15392], bl[15393], bl[15394], bl[15395], bl[15396], bl[15397], bl[15398], bl[15399], bl[15400], bl[15401], bl[15402], bl[15403], bl[15404], bl[15405], bl[15406], bl[15407], bl[15408], bl[15409], bl[15410], bl[15411], bl[15412], bl[15413], bl[15414], bl[15415], bl[15416], bl[15417], bl[15418], bl[15419], bl[15420], bl[15421], bl[15422], bl[15423], bl[15424], bl[15425], bl[15426], bl[15427], bl[15428], bl[15429], bl[15430], bl[15431], bl[15432], bl[15433], bl[15434], bl[15435], bl[15436], bl[15437], bl[15438], bl[15439], bl[15440], bl[15441], bl[15442], bl[15443], bl[15444], bl[15445], bl[15446], bl[15447], bl[15448], bl[15449], bl[15450], bl[15451], bl[15452], bl[15453], bl[15454], bl[15455], bl[16476], bl[16477], bl[16478], bl[16479], bl[16480], bl[16481], bl[16482], bl[16483], bl[16484], bl[16485], bl[16486], bl[16487], bl[16488], bl[16489], bl[16490], bl[16491], bl[16492], bl[16493], bl[16494], bl[16495], bl[16496], bl[16497], bl[16498], bl[16499], bl[16500], bl[16501], bl[16502], bl[16503], bl[16504], bl[16505], bl[16506], bl[16507], bl[16508], bl[16509], bl[16510], bl[16511], bl[16512], bl[16513], bl[16514], bl[16515], bl[16516], bl[16517], bl[16518], bl[16519], bl[16520], bl[16521], bl[16522], bl[16523], bl[16524], bl[16525], bl[16526], bl[16527], bl[16528], bl[16529], bl[16530], bl[16531], bl[16532], bl[16533], bl[16534], bl[16535], bl[16536], bl[16537], bl[16538], bl[16539], bl[16540], bl[16541], bl[16542], bl[16543], bl[16544], bl[16545], bl[16546], bl[16547], bl[16548], bl[16549], bl[16550], bl[16551], bl[16552], bl[16553], bl[16554], bl[16555]}),
        .wl({wl[15456], wl[15457], wl[15458], wl[15459], wl[15460], wl[15461], wl[15462], wl[15463], wl[15464], wl[15465], wl[15466], wl[15467], wl[15468], wl[15469], wl[15470], wl[15471], wl[15472], wl[15473], wl[15474], wl[15475], wl[15476], wl[15477], wl[15478], wl[15479], wl[15480], wl[15481], wl[15482], wl[15483], wl[15484], wl[15485], wl[15486], wl[15487], wl[15488], wl[15489], wl[15490], wl[15491], wl[15492], wl[15493], wl[15494], wl[15495], wl[15496], wl[15497], wl[15498], wl[15499], wl[15500], wl[15501], wl[15502], wl[15503], wl[15504], wl[15505], wl[15506], wl[15507], wl[15508], wl[15509], wl[15510], wl[15511], wl[15512], wl[15513], wl[15514], wl[15515], wl[15516], wl[15517], wl[15518], wl[15519], wl[15520], wl[15521], wl[15522], wl[15523], wl[15524], wl[15525], wl[15526], wl[15527], wl[15528], wl[15529], wl[15530], wl[15531], wl[15532], wl[15533], wl[15534], wl[15535], wl[15536], wl[15537], wl[15538], wl[15539], wl[15540], wl[15541], wl[15542], wl[15543], wl[15544], wl[15545], wl[15546], wl[15547], wl[15548], wl[15549], wl[15550], wl[15551], wl[15552], wl[15553], wl[15554], wl[15555], wl[15556], wl[15557], wl[15558], wl[15559], wl[15560], wl[15561], wl[15562], wl[15563], wl[15564], wl[15565], wl[15566], wl[15567], wl[15568], wl[15569], wl[15570], wl[15571], wl[15572], wl[15573], wl[15574], wl[15575], wl[15576], wl[15577], wl[15578], wl[15579], wl[15580], wl[15581], wl[15582], wl[15583], wl[15584], wl[15585], wl[15586], wl[15587], wl[15588], wl[15589], wl[15590], wl[15591], wl[15592], wl[15593], wl[15594], wl[15595], wl[15596], wl[15597], wl[15598], wl[15599], wl[15600], wl[15601], wl[15602], wl[15603], wl[15604], wl[15605], wl[15606], wl[15607], wl[15608], wl[15609], wl[15610], wl[15611], wl[15612], wl[15613], wl[15614], wl[15615], wl[15616], wl[15617], wl[15618], wl[15619], wl[15620], wl[15621], wl[15622], wl[15623], wl[15624], wl[15625], wl[15626], wl[15627], wl[15628], wl[15629], wl[15630], wl[15631], wl[15632], wl[15633], wl[15634], wl[15635], wl[15636], wl[15637], wl[15638], wl[15639], wl[15640], wl[15641], wl[15642], wl[15643], wl[15644], wl[15645], wl[15646], wl[15647], wl[15648], wl[15649], wl[15650], wl[15651], wl[15652], wl[15653], wl[15654], wl[15655], wl[15656], wl[15657], wl[15658], wl[15659], wl[15660], wl[15661], wl[15662], wl[15663], wl[15664], wl[15665], wl[15666], wl[15667], wl[15668], wl[15669], wl[15670], wl[15671], wl[15672], wl[15673], wl[15674], wl[15675], wl[15676], wl[15677], wl[15678], wl[15679], wl[15680], wl[15681], wl[15682], wl[15683], wl[15684], wl[15685], wl[15686], wl[15687], wl[15688], wl[15689], wl[15690], wl[15691], wl[15692], wl[15693], wl[15694], wl[15695], wl[15696], wl[15697], wl[15698], wl[15699], wl[15700], wl[15701], wl[15702], wl[15703], wl[15704], wl[15705], wl[15706], wl[15707], wl[15708], wl[15709], wl[15710], wl[15711], wl[15712], wl[15713], wl[15714], wl[15715], wl[15716], wl[15717], wl[15718], wl[15719], wl[15720], wl[15721], wl[15722], wl[15723], wl[15724], wl[15725], wl[15726], wl[15727], wl[15728], wl[15729], wl[15730], wl[15731], wl[15732], wl[15733], wl[15734], wl[15735], wl[15736], wl[15737], wl[15738], wl[15739], wl[15740], wl[15741], wl[15742], wl[15743], wl[15744], wl[15745], wl[15746], wl[15747], wl[15748], wl[15749], wl[15750], wl[15751], wl[15752], wl[15753], wl[15754], wl[15755], wl[15756], wl[15757], wl[15758], wl[15759], wl[15760], wl[15761], wl[15762], wl[15763], wl[15764], wl[15765], wl[15766], wl[15767], wl[15768], wl[15769], wl[15770], wl[15771], wl[15772], wl[15773], wl[15774], wl[15775], wl[15776], wl[15777], wl[15778], wl[15779], wl[15780], wl[15781], wl[15782], wl[15783], wl[15784], wl[15785], wl[15786], wl[15787], wl[15788], wl[15789], wl[15790], wl[15791], wl[15792], wl[15793], wl[15794], wl[15795], wl[15796], wl[15797], wl[15798], wl[15799], wl[15800], wl[15801], wl[15802], wl[15803], wl[15804], wl[15805], wl[15806], wl[15807], wl[15808], wl[15809], wl[15810], wl[15811], wl[15812], wl[15813], wl[15814], wl[15815], wl[15816], wl[15817], wl[15818], wl[15819], wl[15820], wl[15821], wl[15822], wl[15823], wl[15824], wl[15825], wl[15826], wl[15827], wl[15828], wl[15829], wl[15830], wl[15831], wl[15832], wl[15833], wl[15834], wl[15835], wl[15836], wl[15837], wl[15838], wl[15839], wl[15840], wl[15841], wl[15842], wl[15843], wl[15844], wl[15845], wl[15846], wl[15847], wl[15848], wl[15849], wl[15850], wl[15851], wl[15852], wl[15853], wl[15854], wl[15855], wl[15856], wl[15857], wl[15858], wl[15859], wl[15860], wl[15861], wl[15862], wl[15863], wl[15864], wl[15865], wl[15866], wl[15867], wl[15868], wl[15869], wl[15870], wl[15871], wl[15872], wl[15873], wl[15874], wl[15875], wl[15876], wl[15877], wl[15878], wl[15879], wl[15880], wl[15881], wl[15882], wl[15883], wl[15884], wl[15885], wl[15886], wl[15887], wl[15888], wl[15889], wl[15890], wl[15891], wl[15892], wl[15893], wl[15894], wl[15895], wl[15896], wl[15897], wl[15898], wl[15899], wl[15900], wl[15901], wl[15902], wl[15903], wl[15904], wl[15905], wl[15906], wl[15907], wl[15908], wl[15909], wl[15910], wl[15911], wl[15912], wl[15913], wl[15914], wl[15915], wl[15916], wl[15917], wl[15918], wl[15919], wl[15920], wl[15921], wl[15922], wl[15923], wl[15924], wl[15925], wl[15926], wl[15927], wl[15928], wl[15929], wl[15930], wl[15931], wl[15932], wl[15933], wl[15934], wl[15935], wl[15936], wl[15937], wl[15938], wl[15939], wl[15940], wl[15941], wl[15942], wl[15943], wl[15944], wl[15945], wl[15946], wl[15947], wl[15948], wl[15949], wl[15950], wl[15951], wl[15952], wl[15953], wl[15954], wl[15955], wl[15956], wl[15957], wl[15958], wl[15959], wl[15960], wl[15961], wl[15962], wl[15963], wl[15964], wl[15965], wl[15966], wl[15967], wl[15968], wl[15969], wl[15970], wl[15971], wl[15972], wl[15973], wl[15974], wl[15975], wl[15976], wl[15977], wl[15978], wl[15979], wl[15980], wl[15981], wl[15982], wl[15983], wl[15984], wl[15985], wl[15986], wl[15987], wl[15988], wl[15989], wl[15990], wl[15991], wl[15992], wl[15993], wl[15994], wl[15995], wl[15996], wl[15997], wl[15998], wl[15999], wl[16000], wl[16001], wl[16002], wl[16003], wl[16004], wl[16005], wl[16006], wl[16007], wl[16008], wl[16009], wl[16010], wl[16011], wl[16012], wl[16013], wl[16014], wl[16015], wl[16016], wl[16017], wl[16018], wl[16019], wl[16020], wl[16021], wl[16022], wl[16023], wl[16024], wl[16025], wl[16026], wl[16027], wl[16028], wl[16029], wl[16030], wl[16031], wl[16032], wl[16033], wl[16034], wl[16035], wl[16036], wl[16037], wl[16038], wl[16039], wl[16040], wl[16041], wl[16042], wl[16043], wl[16044], wl[16045], wl[16046], wl[16047], wl[16048], wl[16049], wl[16050], wl[16051], wl[16052], wl[16053], wl[16054], wl[16055], wl[16056], wl[16057], wl[16058], wl[16059], wl[16060], wl[16061], wl[16062], wl[16063], wl[16064], wl[16065], wl[16066], wl[16067], wl[16068], wl[16069], wl[16070], wl[16071], wl[16072], wl[16073], wl[16074], wl[16075], wl[16076], wl[16077], wl[16078], wl[16079], wl[16080], wl[16081], wl[16082], wl[16083], wl[16084], wl[16085], wl[16086], wl[16087], wl[16088], wl[16089], wl[16090], wl[16091], wl[16092], wl[16093], wl[16094], wl[16095], wl[16096], wl[16097], wl[16098], wl[16099], wl[16100], wl[16101], wl[16102], wl[16103], wl[16104], wl[16105], wl[16106], wl[16107], wl[16108], wl[16109], wl[16110], wl[16111], wl[16112], wl[16113], wl[16114], wl[16115], wl[16116], wl[16117], wl[16118], wl[16119], wl[16120], wl[16121], wl[16122], wl[16123], wl[16124], wl[16125], wl[16126], wl[16127], wl[16128], wl[16129], wl[16130], wl[16131], wl[16132], wl[16133], wl[16134], wl[16135], wl[16136], wl[16137], wl[16138], wl[16139], wl[16140], wl[16141], wl[16142], wl[16143], wl[16144], wl[16145], wl[16146], wl[16147], wl[16148], wl[16149], wl[16150], wl[16151], wl[16152], wl[16153], wl[16154], wl[16155], wl[16156], wl[16157], wl[16158], wl[16159], wl[16160], wl[16161], wl[16162], wl[16163], wl[16164], wl[16165], wl[16166], wl[16167], wl[16168], wl[16169], wl[16170], wl[16171], wl[16172], wl[16173], wl[16174], wl[16175], wl[16176], wl[16177], wl[16178], wl[16179], wl[16180], wl[16181], wl[16182], wl[16183], wl[16184], wl[16185], wl[16186], wl[16187], wl[16188], wl[16189], wl[16190], wl[16191], wl[16192], wl[16193], wl[16194], wl[16195], wl[16196], wl[16197], wl[16198], wl[16199], wl[16200], wl[16201], wl[16202], wl[16203], wl[16204], wl[16205], wl[16206], wl[16207], wl[16208], wl[16209], wl[16210], wl[16211], wl[16212], wl[16213], wl[16214], wl[16215], wl[16216], wl[16217], wl[16218], wl[16219], wl[16220], wl[16221], wl[16222], wl[16223], wl[16224], wl[16225], wl[16226], wl[16227], wl[16228], wl[16229], wl[16230], wl[16231], wl[16232], wl[16233], wl[16234], wl[16235], wl[16236], wl[16237], wl[16238], wl[16239], wl[16240], wl[16241], wl[16242], wl[16243], wl[16244], wl[16245], wl[16246], wl[16247], wl[16248], wl[16249], wl[16250], wl[16251], wl[16252], wl[16253], wl[16254], wl[16255], wl[16256], wl[16257], wl[16258], wl[16259], wl[16260], wl[16261], wl[16262], wl[16263], wl[16264], wl[16265], wl[16266], wl[16267], wl[16268], wl[16269], wl[16270], wl[16271], wl[16272], wl[16273], wl[16274], wl[16275], wl[16276], wl[16277], wl[16278], wl[16279], wl[16280], wl[16281], wl[16282], wl[16283], wl[16284], wl[16285], wl[16286], wl[16287], wl[16288], wl[16289], wl[16290], wl[16291], wl[16292], wl[16293], wl[16294], wl[16295], wl[16296], wl[16297], wl[16298], wl[16299], wl[16300], wl[16301], wl[16302], wl[16303], wl[16304], wl[16305], wl[16306], wl[16307], wl[16308], wl[16309], wl[16310], wl[16311], wl[16312], wl[16313], wl[16314], wl[16315], wl[16316], wl[16317], wl[16318], wl[16319], wl[16320], wl[16321], wl[16322], wl[16323], wl[16324], wl[16325], wl[16326], wl[16327], wl[16328], wl[16329], wl[16330], wl[16331], wl[16332], wl[16333], wl[16334], wl[16335], wl[16336], wl[16337], wl[16338], wl[16339], wl[16340], wl[16341], wl[16342], wl[16343], wl[16344], wl[16345], wl[16346], wl[16347], wl[16348], wl[16349], wl[16350], wl[16351], wl[16352], wl[16353], wl[16354], wl[16355], wl[16356], wl[16357], wl[16358], wl[16359], wl[16360], wl[16361], wl[16362], wl[16363], wl[16364], wl[16365], wl[16366], wl[16367], wl[16368], wl[16369], wl[16370], wl[16371], wl[16372], wl[16373], wl[16374], wl[16375], wl[16376], wl[16377], wl[16378], wl[16379], wl[16380], wl[16381], wl[16382], wl[16383], wl[16384], wl[16385], wl[16386], wl[16387], wl[16388], wl[16389], wl[16390], wl[16391], wl[16392], wl[16393], wl[16394], wl[16395], wl[16396], wl[16397], wl[16398], wl[16399], wl[16400], wl[16401], wl[16402], wl[16403], wl[16404], wl[16405], wl[16406], wl[16407], wl[16408], wl[16409], wl[16410], wl[16411], wl[16412], wl[16413], wl[16414], wl[16415], wl[16416], wl[16417], wl[16418], wl[16419], wl[16420], wl[16421], wl[16422], wl[16423], wl[16424], wl[16425], wl[16426], wl[16427], wl[16428], wl[16429], wl[16430], wl[16431], wl[16432], wl[16433], wl[16434], wl[16435], wl[16436], wl[16437], wl[16438], wl[16439], wl[16440], wl[16441], wl[16442], wl[16443], wl[16444], wl[16445], wl[16446], wl[16447], wl[16448], wl[16449], wl[16450], wl[16451], wl[16452], wl[16453], wl[16454], wl[16455], wl[16456], wl[16457], wl[16458], wl[16459], wl[16460], wl[16461], wl[16462], wl[16463], wl[16464], wl[16465], wl[16466], wl[16467], wl[16468], wl[16469], wl[16470], wl[16471], wl[16472], wl[16473], wl[16474], wl[16475], wl[16556], wl[16557], wl[16558], wl[16559], wl[16560], wl[16561], wl[16562], wl[16563], wl[16564], wl[16565], wl[16566], wl[16567], wl[16568], wl[16569], wl[16570], wl[16571], wl[16572], wl[16573], wl[16574], wl[16575], wl[16576], wl[16577], wl[16578], wl[16579], wl[16580], wl[16581], wl[16582], wl[16583], wl[16584], wl[16585], wl[16586], wl[16587], wl[16588], wl[16589], wl[16590], wl[16591], wl[16592], wl[16593], wl[16594], wl[16595], wl[16596], wl[16597], wl[16598], wl[16599], wl[16600], wl[16601], wl[16602], wl[16603], wl[16604], wl[16605], wl[16606], wl[16607], wl[16608], wl[16609], wl[16610], wl[16611], wl[16612], wl[16613], wl[16614], wl[16615], wl[16616], wl[16617], wl[16618], wl[16619], wl[16620], wl[16621], wl[16622], wl[16623], wl[16624], wl[16625], wl[16626], wl[16627], wl[16628], wl[16629], wl[16630], wl[16631], wl[16632], wl[16633], wl[16634], wl[16635], wl[48], wl[49], wl[50], wl[51], wl[52], wl[53], wl[54], wl[55], wl[15384], wl[15385], wl[15386], wl[15387], wl[15388], wl[15389], wl[15390], wl[15391], wl[15392], wl[15393], wl[15394], wl[15395], wl[15396], wl[15397], wl[15398], wl[15399], wl[15400], wl[15401], wl[15402], wl[15403], wl[15404], wl[15405], wl[15406], wl[15407], wl[15408], wl[15409], wl[15410], wl[15411], wl[15412], wl[15413], wl[15414], wl[15415], wl[15416], wl[15417], wl[15418], wl[15419], wl[15420], wl[15421], wl[15422], wl[15423], wl[15424], wl[15425], wl[15426], wl[15427], wl[15428], wl[15429], wl[15430], wl[15431], wl[15432], wl[15433], wl[15434], wl[15435], wl[15436], wl[15437], wl[15438], wl[15439], wl[15440], wl[15441], wl[15442], wl[15443], wl[15444], wl[15445], wl[15446], wl[15447], wl[15448], wl[15449], wl[15450], wl[15451], wl[15452], wl[15453], wl[15454], wl[15455], wl[16476], wl[16477], wl[16478], wl[16479], wl[16480], wl[16481], wl[16482], wl[16483], wl[16484], wl[16485], wl[16486], wl[16487], wl[16488], wl[16489], wl[16490], wl[16491], wl[16492], wl[16493], wl[16494], wl[16495], wl[16496], wl[16497], wl[16498], wl[16499], wl[16500], wl[16501], wl[16502], wl[16503], wl[16504], wl[16505], wl[16506], wl[16507], wl[16508], wl[16509], wl[16510], wl[16511], wl[16512], wl[16513], wl[16514], wl[16515], wl[16516], wl[16517], wl[16518], wl[16519], wl[16520], wl[16521], wl[16522], wl[16523], wl[16524], wl[16525], wl[16526], wl[16527], wl[16528], wl[16529], wl[16530], wl[16531], wl[16532], wl[16533], wl[16534], wl[16535], wl[16536], wl[16537], wl[16538], wl[16539], wl[16540], wl[16541], wl[16542], wl[16543], wl[16544], wl[16545], wl[16546], wl[16547], wl[16548], wl[16549], wl[16550], wl[16551], wl[16552], wl[16553], wl[16554], wl[16555]})
    );
    top_tile tile_2__5_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_0__4__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_0__4__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_0__4__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_1__3__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_1__3__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_1__3__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_0__3__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_0__3__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_0__3__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_0__3__grid_top_r_in[1]),
        .grid_left_in(grid_clb_1__4__grid_left_in),
        .grid_bottom_in(grid_clb_1__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0:7]),
        .io_bottom_in(grid_io_top_1__5__io_bottom_in),
        .chanx_left_in(sb_0__4__0_chanx_right_out),
        .chanx_left_out(cbx_1__4__0_chanx_left_out),
        .chany_bottom_in(sb_1__1__2_chany_top_out),
        .chany_bottom_out(cby_1__1__3_chany_bottom_out),
        .grid_right_out(grid_clb_2__4__grid_left_in),
        .chanx_right_in_0(cbx_1__4__1_chanx_left_out),
        .chanx_right_out_0(sb_1__4__0_chanx_right_out),
        .grid_right_t_inpad(grid_io_top_2__5__io_bottom_in),
        .grid_right_b_in(sb_1__4__grid_right_b_in),
        .grid_bottom_r_in(sb_1__3__grid_top_r_in),
        .grid_bottom_l_in(sb_1__3__grid_top_l_in),
        .grid_left_b_in(sb_0__4__grid_right_b_in),
        .bl({bl[20488], bl[20489], bl[20490], bl[20491], bl[20492], bl[20493], bl[20494], bl[20495], bl[20496], bl[20497], bl[20498], bl[20499], bl[20500], bl[20501], bl[20502], bl[20503], bl[20504], bl[20505], bl[20506], bl[20507], bl[20508], bl[20509], bl[20510], bl[20511], bl[20512], bl[20513], bl[20514], bl[20515], bl[20516], bl[20517], bl[20518], bl[20519], bl[20520], bl[20521], bl[20522], bl[20523], bl[20524], bl[20525], bl[20526], bl[20527], bl[20528], bl[20529], bl[20530], bl[20531], bl[20532], bl[20533], bl[20534], bl[20535], bl[20536], bl[20537], bl[20538], bl[20539], bl[20540], bl[20541], bl[20542], bl[20543], bl[20544], bl[20545], bl[20546], bl[20547], bl[20548], bl[20549], bl[20550], bl[20551], bl[20552], bl[20553], bl[20554], bl[20555], bl[20556], bl[20557], bl[20558], bl[20559], bl[20560], bl[20561], bl[20562], bl[20563], bl[20564], bl[20565], bl[20566], bl[20567], bl[20568], bl[20569], bl[20570], bl[20571], bl[20572], bl[20573], bl[20574], bl[20575], bl[20576], bl[20577], bl[20578], bl[20579], bl[20580], bl[20581], bl[20582], bl[20583], bl[20584], bl[20585], bl[20586], bl[20587], bl[20588], bl[20589], bl[20590], bl[20591], bl[20592], bl[20593], bl[20594], bl[20595], bl[20596], bl[20597], bl[20598], bl[20599], bl[20600], bl[20601], bl[20602], bl[20603], bl[20604], bl[20605], bl[20606], bl[20607], bl[20608], bl[20609], bl[20610], bl[20611], bl[20612], bl[20613], bl[20614], bl[20615], bl[20616], bl[20617], bl[20618], bl[20619], bl[20620], bl[20621], bl[20622], bl[20623], bl[20624], bl[20625], bl[20626], bl[20627], bl[20628], bl[20629], bl[20630], bl[20631], bl[20632], bl[20633], bl[20634], bl[20635], bl[20636], bl[20637], bl[20638], bl[20639], bl[20640], bl[20641], bl[20642], bl[20643], bl[20644], bl[20645], bl[20646], bl[20647], bl[20648], bl[20649], bl[20650], bl[20651], bl[20652], bl[20653], bl[20654], bl[20655], bl[20656], bl[20657], bl[20658], bl[20659], bl[20660], bl[20661], bl[20662], bl[20663], bl[20664], bl[20665], bl[20666], bl[20667], bl[20668], bl[20669], bl[20670], bl[20671], bl[20672], bl[20673], bl[20674], bl[20675], bl[20676], bl[20677], bl[20678], bl[20679], bl[20680], bl[20681], bl[20682], bl[20683], bl[20684], bl[20685], bl[20686], bl[20687], bl[20688], bl[20689], bl[20690], bl[20691], bl[20692], bl[20693], bl[20694], bl[20695], bl[20696], bl[20697], bl[20698], bl[20699], bl[20700], bl[20701], bl[20702], bl[20703], bl[20704], bl[20705], bl[20706], bl[20707], bl[20708], bl[20709], bl[20710], bl[20711], bl[20712], bl[20713], bl[20714], bl[20715], bl[20716], bl[20717], bl[20718], bl[20719], bl[20720], bl[20721], bl[20722], bl[20723], bl[20724], bl[20725], bl[20726], bl[20727], bl[20728], bl[20729], bl[20730], bl[20731], bl[20732], bl[20733], bl[20734], bl[20735], bl[20736], bl[20737], bl[20738], bl[20739], bl[20740], bl[20741], bl[20742], bl[20743], bl[20744], bl[20745], bl[20746], bl[20747], bl[20748], bl[20749], bl[20750], bl[20751], bl[20752], bl[20753], bl[20754], bl[20755], bl[20756], bl[20757], bl[20758], bl[20759], bl[20760], bl[20761], bl[20762], bl[20763], bl[20764], bl[20765], bl[20766], bl[20767], bl[20768], bl[20769], bl[20770], bl[20771], bl[20772], bl[20773], bl[20774], bl[20775], bl[20776], bl[20777], bl[20778], bl[20779], bl[20780], bl[20781], bl[20782], bl[20783], bl[20784], bl[20785], bl[20786], bl[20787], bl[20788], bl[20789], bl[20790], bl[20791], bl[20792], bl[20793], bl[20794], bl[20795], bl[20796], bl[20797], bl[20798], bl[20799], bl[20800], bl[20801], bl[20802], bl[20803], bl[20804], bl[20805], bl[20806], bl[20807], bl[20808], bl[20809], bl[20810], bl[20811], bl[20812], bl[20813], bl[20814], bl[20815], bl[20816], bl[20817], bl[20818], bl[20819], bl[20820], bl[20821], bl[20822], bl[20823], bl[20824], bl[20825], bl[20826], bl[20827], bl[20828], bl[20829], bl[20830], bl[20831], bl[20832], bl[20833], bl[20834], bl[20835], bl[20836], bl[20837], bl[20838], bl[20839], bl[20840], bl[20841], bl[20842], bl[20843], bl[20844], bl[20845], bl[20846], bl[20847], bl[20848], bl[20849], bl[20850], bl[20851], bl[20852], bl[20853], bl[20854], bl[20855], bl[20856], bl[20857], bl[20858], bl[20859], bl[20860], bl[20861], bl[20862], bl[20863], bl[20864], bl[20865], bl[20866], bl[20867], bl[20868], bl[20869], bl[20870], bl[20871], bl[20872], bl[20873], bl[20874], bl[20875], bl[20876], bl[20877], bl[20878], bl[20879], bl[20880], bl[20881], bl[20882], bl[20883], bl[20884], bl[20885], bl[20886], bl[20887], bl[20888], bl[20889], bl[20890], bl[20891], bl[20892], bl[20893], bl[20894], bl[20895], bl[20896], bl[20897], bl[20898], bl[20899], bl[20900], bl[20901], bl[20902], bl[20903], bl[20904], bl[20905], bl[20906], bl[20907], bl[20908], bl[20909], bl[20910], bl[20911], bl[20912], bl[20913], bl[20914], bl[20915], bl[20916], bl[20917], bl[20918], bl[20919], bl[20920], bl[20921], bl[20922], bl[20923], bl[20924], bl[20925], bl[20926], bl[20927], bl[20928], bl[20929], bl[20930], bl[20931], bl[20932], bl[20933], bl[20934], bl[20935], bl[20936], bl[20937], bl[20938], bl[20939], bl[20940], bl[20941], bl[20942], bl[20943], bl[20944], bl[20945], bl[20946], bl[20947], bl[20948], bl[20949], bl[20950], bl[20951], bl[20952], bl[20953], bl[20954], bl[20955], bl[20956], bl[20957], bl[20958], bl[20959], bl[20960], bl[20961], bl[20962], bl[20963], bl[20964], bl[20965], bl[20966], bl[20967], bl[20968], bl[20969], bl[20970], bl[20971], bl[20972], bl[20973], bl[20974], bl[20975], bl[20976], bl[20977], bl[20978], bl[20979], bl[20980], bl[20981], bl[20982], bl[20983], bl[20984], bl[20985], bl[20986], bl[20987], bl[20988], bl[20989], bl[20990], bl[20991], bl[20992], bl[20993], bl[20994], bl[20995], bl[20996], bl[20997], bl[20998], bl[20999], bl[21000], bl[21001], bl[21002], bl[21003], bl[21004], bl[21005], bl[21006], bl[21007], bl[21008], bl[21009], bl[21010], bl[21011], bl[21012], bl[21013], bl[21014], bl[21015], bl[21016], bl[21017], bl[21018], bl[21019], bl[21020], bl[21021], bl[21022], bl[21023], bl[21024], bl[21025], bl[21026], bl[21027], bl[21028], bl[21029], bl[21030], bl[21031], bl[21032], bl[21033], bl[21034], bl[21035], bl[21036], bl[21037], bl[21038], bl[21039], bl[21040], bl[21041], bl[21042], bl[21043], bl[21044], bl[21045], bl[21046], bl[21047], bl[21048], bl[21049], bl[21050], bl[21051], bl[21052], bl[21053], bl[21054], bl[21055], bl[21056], bl[21057], bl[21058], bl[21059], bl[21060], bl[21061], bl[21062], bl[21063], bl[21064], bl[21065], bl[21066], bl[21067], bl[21068], bl[21069], bl[21070], bl[21071], bl[21072], bl[21073], bl[21074], bl[21075], bl[21076], bl[21077], bl[21078], bl[21079], bl[21080], bl[21081], bl[21082], bl[21083], bl[21084], bl[21085], bl[21086], bl[21087], bl[21088], bl[21089], bl[21090], bl[21091], bl[21092], bl[21093], bl[21094], bl[21095], bl[21096], bl[21097], bl[21098], bl[21099], bl[21100], bl[21101], bl[21102], bl[21103], bl[21104], bl[21105], bl[21106], bl[21107], bl[21108], bl[21109], bl[21110], bl[21111], bl[21112], bl[21113], bl[21114], bl[21115], bl[21116], bl[21117], bl[21118], bl[21119], bl[21120], bl[21121], bl[21122], bl[21123], bl[21124], bl[21125], bl[21126], bl[21127], bl[21128], bl[21129], bl[21130], bl[21131], bl[21132], bl[21133], bl[21134], bl[21135], bl[21136], bl[21137], bl[21138], bl[21139], bl[21140], bl[21141], bl[21142], bl[21143], bl[21144], bl[21145], bl[21146], bl[21147], bl[21148], bl[21149], bl[21150], bl[21151], bl[21152], bl[21153], bl[21154], bl[21155], bl[21156], bl[21157], bl[21158], bl[21159], bl[21160], bl[21161], bl[21162], bl[21163], bl[21164], bl[21165], bl[21166], bl[21167], bl[21168], bl[21169], bl[21170], bl[21171], bl[21172], bl[21173], bl[21174], bl[21175], bl[21176], bl[21177], bl[21178], bl[21179], bl[21180], bl[21181], bl[21182], bl[21183], bl[21184], bl[21185], bl[21186], bl[21187], bl[21188], bl[21189], bl[21190], bl[21191], bl[21192], bl[21193], bl[21194], bl[21195], bl[21196], bl[21197], bl[21198], bl[21199], bl[21200], bl[21201], bl[21202], bl[21203], bl[21204], bl[21205], bl[21206], bl[21207], bl[21208], bl[21209], bl[21210], bl[21211], bl[21212], bl[21213], bl[21214], bl[21215], bl[21216], bl[21217], bl[21218], bl[21219], bl[21220], bl[21221], bl[21222], bl[21223], bl[21224], bl[21225], bl[21226], bl[21227], bl[21228], bl[21229], bl[21230], bl[21231], bl[21232], bl[21233], bl[21234], bl[21235], bl[21236], bl[21237], bl[21238], bl[21239], bl[21240], bl[21241], bl[21242], bl[21243], bl[21244], bl[21245], bl[21246], bl[21247], bl[21248], bl[21249], bl[21250], bl[21251], bl[21252], bl[21253], bl[21254], bl[21255], bl[21256], bl[21257], bl[21258], bl[21259], bl[21260], bl[21261], bl[21262], bl[21263], bl[21264], bl[21265], bl[21266], bl[21267], bl[21268], bl[21269], bl[21270], bl[21271], bl[21272], bl[21273], bl[21274], bl[21275], bl[21276], bl[21277], bl[21278], bl[21279], bl[21280], bl[21281], bl[21282], bl[21283], bl[21284], bl[21285], bl[21286], bl[21287], bl[21288], bl[21289], bl[21290], bl[21291], bl[21292], bl[21293], bl[21294], bl[21295], bl[21296], bl[21297], bl[21298], bl[21299], bl[21300], bl[21301], bl[21302], bl[21303], bl[21304], bl[21305], bl[21306], bl[21307], bl[21308], bl[21309], bl[21310], bl[21311], bl[21312], bl[21313], bl[21314], bl[21315], bl[21316], bl[21317], bl[21318], bl[21319], bl[21320], bl[21321], bl[21322], bl[21323], bl[21324], bl[21325], bl[21326], bl[21327], bl[21328], bl[21329], bl[21330], bl[21331], bl[21332], bl[21333], bl[21334], bl[21335], bl[21336], bl[21337], bl[21338], bl[21339], bl[21340], bl[21341], bl[21342], bl[21343], bl[21344], bl[21345], bl[21346], bl[21347], bl[21348], bl[21349], bl[21350], bl[21351], bl[21352], bl[21353], bl[21354], bl[21355], bl[21356], bl[21357], bl[21358], bl[21359], bl[21360], bl[21361], bl[21362], bl[21363], bl[21364], bl[21365], bl[21366], bl[21367], bl[21368], bl[21369], bl[21370], bl[21371], bl[21372], bl[21373], bl[21374], bl[21375], bl[21376], bl[21377], bl[21378], bl[21379], bl[21380], bl[21381], bl[21382], bl[21383], bl[21384], bl[21385], bl[21386], bl[21387], bl[21388], bl[21389], bl[21390], bl[21391], bl[21392], bl[21393], bl[21394], bl[21395], bl[21396], bl[21397], bl[21398], bl[21399], bl[21400], bl[21401], bl[21402], bl[21403], bl[21404], bl[21405], bl[21406], bl[21407], bl[21408], bl[21409], bl[21410], bl[21411], bl[21412], bl[21413], bl[21414], bl[21415], bl[21416], bl[21417], bl[21418], bl[21419], bl[21420], bl[21421], bl[21422], bl[21423], bl[21424], bl[21425], bl[21426], bl[21427], bl[21428], bl[21429], bl[21430], bl[21431], bl[21432], bl[21433], bl[21434], bl[21435], bl[21436], bl[21437], bl[21438], bl[21439], bl[21440], bl[21441], bl[21442], bl[21443], bl[21444], bl[21445], bl[21446], bl[21447], bl[21448], bl[21449], bl[21450], bl[21451], bl[21452], bl[21453], bl[21454], bl[21455], bl[21456], bl[21457], bl[21458], bl[21459], bl[21460], bl[21461], bl[21462], bl[21463], bl[21464], bl[21465], bl[21466], bl[21467], bl[21468], bl[21469], bl[21470], bl[21471], bl[21472], bl[21473], bl[21474], bl[21475], bl[21476], bl[21477], bl[21478], bl[21479], bl[21480], bl[21481], bl[21482], bl[21483], bl[21484], bl[21485], bl[21486], bl[21487], bl[21488], bl[21489], bl[21490], bl[21491], bl[21492], bl[21493], bl[21494], bl[21495], bl[21496], bl[21497], bl[21498], bl[21499], bl[21500], bl[21501], bl[21502], bl[21503], bl[21504], bl[21505], bl[21506], bl[21507], bl[696], bl[697], bl[698], bl[699], bl[700], bl[701], bl[702], bl[703], bl[624], bl[625], bl[626], bl[627], bl[628], bl[629], bl[630], bl[631], bl[632], bl[633], bl[634], bl[635], bl[636], bl[637], bl[638], bl[639], bl[640], bl[641], bl[642], bl[643], bl[644], bl[645], bl[646], bl[647], bl[648], bl[649], bl[650], bl[651], bl[652], bl[653], bl[654], bl[655], bl[656], bl[657], bl[658], bl[659], bl[660], bl[661], bl[662], bl[663], bl[664], bl[665], bl[666], bl[667], bl[668], bl[669], bl[670], bl[671], bl[672], bl[673], bl[674], bl[675], bl[676], bl[677], bl[678], bl[679], bl[680], bl[681], bl[682], bl[683], bl[684], bl[685], bl[686], bl[687], bl[688], bl[689], bl[690], bl[691], bl[692], bl[693], bl[694], bl[695], bl[20408], bl[20409], bl[20410], bl[20411], bl[20412], bl[20413], bl[20414], bl[20415], bl[20416], bl[20417], bl[20418], bl[20419], bl[20420], bl[20421], bl[20422], bl[20423], bl[20424], bl[20425], bl[20426], bl[20427], bl[20428], bl[20429], bl[20430], bl[20431], bl[20432], bl[20433], bl[20434], bl[20435], bl[20436], bl[20437], bl[20438], bl[20439], bl[20440], bl[20441], bl[20442], bl[20443], bl[20444], bl[20445], bl[20446], bl[20447], bl[20448], bl[20449], bl[20450], bl[20451], bl[20452], bl[20453], bl[20454], bl[20455], bl[20456], bl[20457], bl[20458], bl[20459], bl[20460], bl[20461], bl[20462], bl[20463], bl[20464], bl[20465], bl[20466], bl[20467], bl[20468], bl[20469], bl[20470], bl[20471], bl[20472], bl[20473], bl[20474], bl[20475], bl[20476], bl[20477], bl[20478], bl[20479], bl[20480], bl[20481], bl[20482], bl[20483], bl[20484], bl[20485], bl[20486], bl[20487], bl[544], bl[545], bl[546], bl[547], bl[548], bl[549], bl[550], bl[551], bl[552], bl[553], bl[554], bl[555], bl[556], bl[557], bl[558], bl[559], bl[560], bl[561], bl[562], bl[563], bl[564], bl[565], bl[566], bl[567], bl[568], bl[569], bl[570], bl[571], bl[572], bl[573], bl[574], bl[575], bl[576], bl[577], bl[578], bl[579], bl[580], bl[581], bl[582], bl[583], bl[584], bl[585], bl[586], bl[587], bl[588], bl[589], bl[590], bl[591], bl[592], bl[593], bl[594], bl[595], bl[596], bl[597], bl[598], bl[599], bl[600], bl[601], bl[602], bl[603], bl[604], bl[605], bl[606], bl[607], bl[608], bl[609], bl[610], bl[611], bl[612], bl[613], bl[614], bl[615], bl[616], bl[617], bl[618], bl[619], bl[620], bl[621], bl[622], bl[623]}),
        .wl({wl[20488], wl[20489], wl[20490], wl[20491], wl[20492], wl[20493], wl[20494], wl[20495], wl[20496], wl[20497], wl[20498], wl[20499], wl[20500], wl[20501], wl[20502], wl[20503], wl[20504], wl[20505], wl[20506], wl[20507], wl[20508], wl[20509], wl[20510], wl[20511], wl[20512], wl[20513], wl[20514], wl[20515], wl[20516], wl[20517], wl[20518], wl[20519], wl[20520], wl[20521], wl[20522], wl[20523], wl[20524], wl[20525], wl[20526], wl[20527], wl[20528], wl[20529], wl[20530], wl[20531], wl[20532], wl[20533], wl[20534], wl[20535], wl[20536], wl[20537], wl[20538], wl[20539], wl[20540], wl[20541], wl[20542], wl[20543], wl[20544], wl[20545], wl[20546], wl[20547], wl[20548], wl[20549], wl[20550], wl[20551], wl[20552], wl[20553], wl[20554], wl[20555], wl[20556], wl[20557], wl[20558], wl[20559], wl[20560], wl[20561], wl[20562], wl[20563], wl[20564], wl[20565], wl[20566], wl[20567], wl[20568], wl[20569], wl[20570], wl[20571], wl[20572], wl[20573], wl[20574], wl[20575], wl[20576], wl[20577], wl[20578], wl[20579], wl[20580], wl[20581], wl[20582], wl[20583], wl[20584], wl[20585], wl[20586], wl[20587], wl[20588], wl[20589], wl[20590], wl[20591], wl[20592], wl[20593], wl[20594], wl[20595], wl[20596], wl[20597], wl[20598], wl[20599], wl[20600], wl[20601], wl[20602], wl[20603], wl[20604], wl[20605], wl[20606], wl[20607], wl[20608], wl[20609], wl[20610], wl[20611], wl[20612], wl[20613], wl[20614], wl[20615], wl[20616], wl[20617], wl[20618], wl[20619], wl[20620], wl[20621], wl[20622], wl[20623], wl[20624], wl[20625], wl[20626], wl[20627], wl[20628], wl[20629], wl[20630], wl[20631], wl[20632], wl[20633], wl[20634], wl[20635], wl[20636], wl[20637], wl[20638], wl[20639], wl[20640], wl[20641], wl[20642], wl[20643], wl[20644], wl[20645], wl[20646], wl[20647], wl[20648], wl[20649], wl[20650], wl[20651], wl[20652], wl[20653], wl[20654], wl[20655], wl[20656], wl[20657], wl[20658], wl[20659], wl[20660], wl[20661], wl[20662], wl[20663], wl[20664], wl[20665], wl[20666], wl[20667], wl[20668], wl[20669], wl[20670], wl[20671], wl[20672], wl[20673], wl[20674], wl[20675], wl[20676], wl[20677], wl[20678], wl[20679], wl[20680], wl[20681], wl[20682], wl[20683], wl[20684], wl[20685], wl[20686], wl[20687], wl[20688], wl[20689], wl[20690], wl[20691], wl[20692], wl[20693], wl[20694], wl[20695], wl[20696], wl[20697], wl[20698], wl[20699], wl[20700], wl[20701], wl[20702], wl[20703], wl[20704], wl[20705], wl[20706], wl[20707], wl[20708], wl[20709], wl[20710], wl[20711], wl[20712], wl[20713], wl[20714], wl[20715], wl[20716], wl[20717], wl[20718], wl[20719], wl[20720], wl[20721], wl[20722], wl[20723], wl[20724], wl[20725], wl[20726], wl[20727], wl[20728], wl[20729], wl[20730], wl[20731], wl[20732], wl[20733], wl[20734], wl[20735], wl[20736], wl[20737], wl[20738], wl[20739], wl[20740], wl[20741], wl[20742], wl[20743], wl[20744], wl[20745], wl[20746], wl[20747], wl[20748], wl[20749], wl[20750], wl[20751], wl[20752], wl[20753], wl[20754], wl[20755], wl[20756], wl[20757], wl[20758], wl[20759], wl[20760], wl[20761], wl[20762], wl[20763], wl[20764], wl[20765], wl[20766], wl[20767], wl[20768], wl[20769], wl[20770], wl[20771], wl[20772], wl[20773], wl[20774], wl[20775], wl[20776], wl[20777], wl[20778], wl[20779], wl[20780], wl[20781], wl[20782], wl[20783], wl[20784], wl[20785], wl[20786], wl[20787], wl[20788], wl[20789], wl[20790], wl[20791], wl[20792], wl[20793], wl[20794], wl[20795], wl[20796], wl[20797], wl[20798], wl[20799], wl[20800], wl[20801], wl[20802], wl[20803], wl[20804], wl[20805], wl[20806], wl[20807], wl[20808], wl[20809], wl[20810], wl[20811], wl[20812], wl[20813], wl[20814], wl[20815], wl[20816], wl[20817], wl[20818], wl[20819], wl[20820], wl[20821], wl[20822], wl[20823], wl[20824], wl[20825], wl[20826], wl[20827], wl[20828], wl[20829], wl[20830], wl[20831], wl[20832], wl[20833], wl[20834], wl[20835], wl[20836], wl[20837], wl[20838], wl[20839], wl[20840], wl[20841], wl[20842], wl[20843], wl[20844], wl[20845], wl[20846], wl[20847], wl[20848], wl[20849], wl[20850], wl[20851], wl[20852], wl[20853], wl[20854], wl[20855], wl[20856], wl[20857], wl[20858], wl[20859], wl[20860], wl[20861], wl[20862], wl[20863], wl[20864], wl[20865], wl[20866], wl[20867], wl[20868], wl[20869], wl[20870], wl[20871], wl[20872], wl[20873], wl[20874], wl[20875], wl[20876], wl[20877], wl[20878], wl[20879], wl[20880], wl[20881], wl[20882], wl[20883], wl[20884], wl[20885], wl[20886], wl[20887], wl[20888], wl[20889], wl[20890], wl[20891], wl[20892], wl[20893], wl[20894], wl[20895], wl[20896], wl[20897], wl[20898], wl[20899], wl[20900], wl[20901], wl[20902], wl[20903], wl[20904], wl[20905], wl[20906], wl[20907], wl[20908], wl[20909], wl[20910], wl[20911], wl[20912], wl[20913], wl[20914], wl[20915], wl[20916], wl[20917], wl[20918], wl[20919], wl[20920], wl[20921], wl[20922], wl[20923], wl[20924], wl[20925], wl[20926], wl[20927], wl[20928], wl[20929], wl[20930], wl[20931], wl[20932], wl[20933], wl[20934], wl[20935], wl[20936], wl[20937], wl[20938], wl[20939], wl[20940], wl[20941], wl[20942], wl[20943], wl[20944], wl[20945], wl[20946], wl[20947], wl[20948], wl[20949], wl[20950], wl[20951], wl[20952], wl[20953], wl[20954], wl[20955], wl[20956], wl[20957], wl[20958], wl[20959], wl[20960], wl[20961], wl[20962], wl[20963], wl[20964], wl[20965], wl[20966], wl[20967], wl[20968], wl[20969], wl[20970], wl[20971], wl[20972], wl[20973], wl[20974], wl[20975], wl[20976], wl[20977], wl[20978], wl[20979], wl[20980], wl[20981], wl[20982], wl[20983], wl[20984], wl[20985], wl[20986], wl[20987], wl[20988], wl[20989], wl[20990], wl[20991], wl[20992], wl[20993], wl[20994], wl[20995], wl[20996], wl[20997], wl[20998], wl[20999], wl[21000], wl[21001], wl[21002], wl[21003], wl[21004], wl[21005], wl[21006], wl[21007], wl[21008], wl[21009], wl[21010], wl[21011], wl[21012], wl[21013], wl[21014], wl[21015], wl[21016], wl[21017], wl[21018], wl[21019], wl[21020], wl[21021], wl[21022], wl[21023], wl[21024], wl[21025], wl[21026], wl[21027], wl[21028], wl[21029], wl[21030], wl[21031], wl[21032], wl[21033], wl[21034], wl[21035], wl[21036], wl[21037], wl[21038], wl[21039], wl[21040], wl[21041], wl[21042], wl[21043], wl[21044], wl[21045], wl[21046], wl[21047], wl[21048], wl[21049], wl[21050], wl[21051], wl[21052], wl[21053], wl[21054], wl[21055], wl[21056], wl[21057], wl[21058], wl[21059], wl[21060], wl[21061], wl[21062], wl[21063], wl[21064], wl[21065], wl[21066], wl[21067], wl[21068], wl[21069], wl[21070], wl[21071], wl[21072], wl[21073], wl[21074], wl[21075], wl[21076], wl[21077], wl[21078], wl[21079], wl[21080], wl[21081], wl[21082], wl[21083], wl[21084], wl[21085], wl[21086], wl[21087], wl[21088], wl[21089], wl[21090], wl[21091], wl[21092], wl[21093], wl[21094], wl[21095], wl[21096], wl[21097], wl[21098], wl[21099], wl[21100], wl[21101], wl[21102], wl[21103], wl[21104], wl[21105], wl[21106], wl[21107], wl[21108], wl[21109], wl[21110], wl[21111], wl[21112], wl[21113], wl[21114], wl[21115], wl[21116], wl[21117], wl[21118], wl[21119], wl[21120], wl[21121], wl[21122], wl[21123], wl[21124], wl[21125], wl[21126], wl[21127], wl[21128], wl[21129], wl[21130], wl[21131], wl[21132], wl[21133], wl[21134], wl[21135], wl[21136], wl[21137], wl[21138], wl[21139], wl[21140], wl[21141], wl[21142], wl[21143], wl[21144], wl[21145], wl[21146], wl[21147], wl[21148], wl[21149], wl[21150], wl[21151], wl[21152], wl[21153], wl[21154], wl[21155], wl[21156], wl[21157], wl[21158], wl[21159], wl[21160], wl[21161], wl[21162], wl[21163], wl[21164], wl[21165], wl[21166], wl[21167], wl[21168], wl[21169], wl[21170], wl[21171], wl[21172], wl[21173], wl[21174], wl[21175], wl[21176], wl[21177], wl[21178], wl[21179], wl[21180], wl[21181], wl[21182], wl[21183], wl[21184], wl[21185], wl[21186], wl[21187], wl[21188], wl[21189], wl[21190], wl[21191], wl[21192], wl[21193], wl[21194], wl[21195], wl[21196], wl[21197], wl[21198], wl[21199], wl[21200], wl[21201], wl[21202], wl[21203], wl[21204], wl[21205], wl[21206], wl[21207], wl[21208], wl[21209], wl[21210], wl[21211], wl[21212], wl[21213], wl[21214], wl[21215], wl[21216], wl[21217], wl[21218], wl[21219], wl[21220], wl[21221], wl[21222], wl[21223], wl[21224], wl[21225], wl[21226], wl[21227], wl[21228], wl[21229], wl[21230], wl[21231], wl[21232], wl[21233], wl[21234], wl[21235], wl[21236], wl[21237], wl[21238], wl[21239], wl[21240], wl[21241], wl[21242], wl[21243], wl[21244], wl[21245], wl[21246], wl[21247], wl[21248], wl[21249], wl[21250], wl[21251], wl[21252], wl[21253], wl[21254], wl[21255], wl[21256], wl[21257], wl[21258], wl[21259], wl[21260], wl[21261], wl[21262], wl[21263], wl[21264], wl[21265], wl[21266], wl[21267], wl[21268], wl[21269], wl[21270], wl[21271], wl[21272], wl[21273], wl[21274], wl[21275], wl[21276], wl[21277], wl[21278], wl[21279], wl[21280], wl[21281], wl[21282], wl[21283], wl[21284], wl[21285], wl[21286], wl[21287], wl[21288], wl[21289], wl[21290], wl[21291], wl[21292], wl[21293], wl[21294], wl[21295], wl[21296], wl[21297], wl[21298], wl[21299], wl[21300], wl[21301], wl[21302], wl[21303], wl[21304], wl[21305], wl[21306], wl[21307], wl[21308], wl[21309], wl[21310], wl[21311], wl[21312], wl[21313], wl[21314], wl[21315], wl[21316], wl[21317], wl[21318], wl[21319], wl[21320], wl[21321], wl[21322], wl[21323], wl[21324], wl[21325], wl[21326], wl[21327], wl[21328], wl[21329], wl[21330], wl[21331], wl[21332], wl[21333], wl[21334], wl[21335], wl[21336], wl[21337], wl[21338], wl[21339], wl[21340], wl[21341], wl[21342], wl[21343], wl[21344], wl[21345], wl[21346], wl[21347], wl[21348], wl[21349], wl[21350], wl[21351], wl[21352], wl[21353], wl[21354], wl[21355], wl[21356], wl[21357], wl[21358], wl[21359], wl[21360], wl[21361], wl[21362], wl[21363], wl[21364], wl[21365], wl[21366], wl[21367], wl[21368], wl[21369], wl[21370], wl[21371], wl[21372], wl[21373], wl[21374], wl[21375], wl[21376], wl[21377], wl[21378], wl[21379], wl[21380], wl[21381], wl[21382], wl[21383], wl[21384], wl[21385], wl[21386], wl[21387], wl[21388], wl[21389], wl[21390], wl[21391], wl[21392], wl[21393], wl[21394], wl[21395], wl[21396], wl[21397], wl[21398], wl[21399], wl[21400], wl[21401], wl[21402], wl[21403], wl[21404], wl[21405], wl[21406], wl[21407], wl[21408], wl[21409], wl[21410], wl[21411], wl[21412], wl[21413], wl[21414], wl[21415], wl[21416], wl[21417], wl[21418], wl[21419], wl[21420], wl[21421], wl[21422], wl[21423], wl[21424], wl[21425], wl[21426], wl[21427], wl[21428], wl[21429], wl[21430], wl[21431], wl[21432], wl[21433], wl[21434], wl[21435], wl[21436], wl[21437], wl[21438], wl[21439], wl[21440], wl[21441], wl[21442], wl[21443], wl[21444], wl[21445], wl[21446], wl[21447], wl[21448], wl[21449], wl[21450], wl[21451], wl[21452], wl[21453], wl[21454], wl[21455], wl[21456], wl[21457], wl[21458], wl[21459], wl[21460], wl[21461], wl[21462], wl[21463], wl[21464], wl[21465], wl[21466], wl[21467], wl[21468], wl[21469], wl[21470], wl[21471], wl[21472], wl[21473], wl[21474], wl[21475], wl[21476], wl[21477], wl[21478], wl[21479], wl[21480], wl[21481], wl[21482], wl[21483], wl[21484], wl[21485], wl[21486], wl[21487], wl[21488], wl[21489], wl[21490], wl[21491], wl[21492], wl[21493], wl[21494], wl[21495], wl[21496], wl[21497], wl[21498], wl[21499], wl[21500], wl[21501], wl[21502], wl[21503], wl[21504], wl[21505], wl[21506], wl[21507], wl[696], wl[697], wl[698], wl[699], wl[700], wl[701], wl[702], wl[703], wl[624], wl[625], wl[626], wl[627], wl[628], wl[629], wl[630], wl[631], wl[632], wl[633], wl[634], wl[635], wl[636], wl[637], wl[638], wl[639], wl[640], wl[641], wl[642], wl[643], wl[644], wl[645], wl[646], wl[647], wl[648], wl[649], wl[650], wl[651], wl[652], wl[653], wl[654], wl[655], wl[656], wl[657], wl[658], wl[659], wl[660], wl[661], wl[662], wl[663], wl[664], wl[665], wl[666], wl[667], wl[668], wl[669], wl[670], wl[671], wl[672], wl[673], wl[674], wl[675], wl[676], wl[677], wl[678], wl[679], wl[680], wl[681], wl[682], wl[683], wl[684], wl[685], wl[686], wl[687], wl[688], wl[689], wl[690], wl[691], wl[692], wl[693], wl[694], wl[695], wl[20408], wl[20409], wl[20410], wl[20411], wl[20412], wl[20413], wl[20414], wl[20415], wl[20416], wl[20417], wl[20418], wl[20419], wl[20420], wl[20421], wl[20422], wl[20423], wl[20424], wl[20425], wl[20426], wl[20427], wl[20428], wl[20429], wl[20430], wl[20431], wl[20432], wl[20433], wl[20434], wl[20435], wl[20436], wl[20437], wl[20438], wl[20439], wl[20440], wl[20441], wl[20442], wl[20443], wl[20444], wl[20445], wl[20446], wl[20447], wl[20448], wl[20449], wl[20450], wl[20451], wl[20452], wl[20453], wl[20454], wl[20455], wl[20456], wl[20457], wl[20458], wl[20459], wl[20460], wl[20461], wl[20462], wl[20463], wl[20464], wl[20465], wl[20466], wl[20467], wl[20468], wl[20469], wl[20470], wl[20471], wl[20472], wl[20473], wl[20474], wl[20475], wl[20476], wl[20477], wl[20478], wl[20479], wl[20480], wl[20481], wl[20482], wl[20483], wl[20484], wl[20485], wl[20486], wl[20487], wl[544], wl[545], wl[546], wl[547], wl[548], wl[549], wl[550], wl[551], wl[552], wl[553], wl[554], wl[555], wl[556], wl[557], wl[558], wl[559], wl[560], wl[561], wl[562], wl[563], wl[564], wl[565], wl[566], wl[567], wl[568], wl[569], wl[570], wl[571], wl[572], wl[573], wl[574], wl[575], wl[576], wl[577], wl[578], wl[579], wl[580], wl[581], wl[582], wl[583], wl[584], wl[585], wl[586], wl[587], wl[588], wl[589], wl[590], wl[591], wl[592], wl[593], wl[594], wl[595], wl[596], wl[597], wl[598], wl[599], wl[600], wl[601], wl[602], wl[603], wl[604], wl[605], wl[606], wl[607], wl[608], wl[609], wl[610], wl[611], wl[612], wl[613], wl[614], wl[615], wl[616], wl[617], wl[618], wl[619], wl[620], wl[621], wl[622], wl[623]})
    );
    top_tile tile_3__5_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_1__4__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_1__4__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_1__4__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_2__3__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_2__3__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_2__3__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_1__3__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_1__3__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_1__3__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_1__3__grid_top_r_in[1]),
        .grid_left_in(grid_clb_2__4__grid_left_in),
        .grid_bottom_in(grid_clb_2__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[8:15]),
        .io_bottom_in(grid_io_top_2__5__io_bottom_in),
        .chanx_left_in(sb_1__4__0_chanx_right_out),
        .chanx_left_out(cbx_1__4__1_chanx_left_out),
        .chany_bottom_in(sb_1__1__5_chany_top_out),
        .chany_bottom_out(cby_1__1__7_chany_bottom_out),
        .grid_right_out(grid_clb_3__4__grid_left_in),
        .chanx_right_in_0(cbx_1__4__2_chanx_left_out),
        .chanx_right_out_0(sb_1__4__1_chanx_right_out),
        .grid_right_t_inpad(grid_io_top_3__5__io_bottom_in),
        .grid_right_b_in(sb_2__4__grid_right_b_in),
        .grid_bottom_r_in(sb_2__3__grid_top_r_in),
        .grid_bottom_l_in(sb_2__3__grid_top_l_in),
        .grid_left_b_in(sb_1__4__grid_right_b_in),
        .bl({bl[19228], bl[19229], bl[19230], bl[19231], bl[19232], bl[19233], bl[19234], bl[19235], bl[19236], bl[19237], bl[19238], bl[19239], bl[19240], bl[19241], bl[19242], bl[19243], bl[19244], bl[19245], bl[19246], bl[19247], bl[19248], bl[19249], bl[19250], bl[19251], bl[19252], bl[19253], bl[19254], bl[19255], bl[19256], bl[19257], bl[19258], bl[19259], bl[19260], bl[19261], bl[19262], bl[19263], bl[19264], bl[19265], bl[19266], bl[19267], bl[19268], bl[19269], bl[19270], bl[19271], bl[19272], bl[19273], bl[19274], bl[19275], bl[19276], bl[19277], bl[19278], bl[19279], bl[19280], bl[19281], bl[19282], bl[19283], bl[19284], bl[19285], bl[19286], bl[19287], bl[19288], bl[19289], bl[19290], bl[19291], bl[19292], bl[19293], bl[19294], bl[19295], bl[19296], bl[19297], bl[19298], bl[19299], bl[19300], bl[19301], bl[19302], bl[19303], bl[19304], bl[19305], bl[19306], bl[19307], bl[19308], bl[19309], bl[19310], bl[19311], bl[19312], bl[19313], bl[19314], bl[19315], bl[19316], bl[19317], bl[19318], bl[19319], bl[19320], bl[19321], bl[19322], bl[19323], bl[19324], bl[19325], bl[19326], bl[19327], bl[19328], bl[19329], bl[19330], bl[19331], bl[19332], bl[19333], bl[19334], bl[19335], bl[19336], bl[19337], bl[19338], bl[19339], bl[19340], bl[19341], bl[19342], bl[19343], bl[19344], bl[19345], bl[19346], bl[19347], bl[19348], bl[19349], bl[19350], bl[19351], bl[19352], bl[19353], bl[19354], bl[19355], bl[19356], bl[19357], bl[19358], bl[19359], bl[19360], bl[19361], bl[19362], bl[19363], bl[19364], bl[19365], bl[19366], bl[19367], bl[19368], bl[19369], bl[19370], bl[19371], bl[19372], bl[19373], bl[19374], bl[19375], bl[19376], bl[19377], bl[19378], bl[19379], bl[19380], bl[19381], bl[19382], bl[19383], bl[19384], bl[19385], bl[19386], bl[19387], bl[19388], bl[19389], bl[19390], bl[19391], bl[19392], bl[19393], bl[19394], bl[19395], bl[19396], bl[19397], bl[19398], bl[19399], bl[19400], bl[19401], bl[19402], bl[19403], bl[19404], bl[19405], bl[19406], bl[19407], bl[19408], bl[19409], bl[19410], bl[19411], bl[19412], bl[19413], bl[19414], bl[19415], bl[19416], bl[19417], bl[19418], bl[19419], bl[19420], bl[19421], bl[19422], bl[19423], bl[19424], bl[19425], bl[19426], bl[19427], bl[19428], bl[19429], bl[19430], bl[19431], bl[19432], bl[19433], bl[19434], bl[19435], bl[19436], bl[19437], bl[19438], bl[19439], bl[19440], bl[19441], bl[19442], bl[19443], bl[19444], bl[19445], bl[19446], bl[19447], bl[19448], bl[19449], bl[19450], bl[19451], bl[19452], bl[19453], bl[19454], bl[19455], bl[19456], bl[19457], bl[19458], bl[19459], bl[19460], bl[19461], bl[19462], bl[19463], bl[19464], bl[19465], bl[19466], bl[19467], bl[19468], bl[19469], bl[19470], bl[19471], bl[19472], bl[19473], bl[19474], bl[19475], bl[19476], bl[19477], bl[19478], bl[19479], bl[19480], bl[19481], bl[19482], bl[19483], bl[19484], bl[19485], bl[19486], bl[19487], bl[19488], bl[19489], bl[19490], bl[19491], bl[19492], bl[19493], bl[19494], bl[19495], bl[19496], bl[19497], bl[19498], bl[19499], bl[19500], bl[19501], bl[19502], bl[19503], bl[19504], bl[19505], bl[19506], bl[19507], bl[19508], bl[19509], bl[19510], bl[19511], bl[19512], bl[19513], bl[19514], bl[19515], bl[19516], bl[19517], bl[19518], bl[19519], bl[19520], bl[19521], bl[19522], bl[19523], bl[19524], bl[19525], bl[19526], bl[19527], bl[19528], bl[19529], bl[19530], bl[19531], bl[19532], bl[19533], bl[19534], bl[19535], bl[19536], bl[19537], bl[19538], bl[19539], bl[19540], bl[19541], bl[19542], bl[19543], bl[19544], bl[19545], bl[19546], bl[19547], bl[19548], bl[19549], bl[19550], bl[19551], bl[19552], bl[19553], bl[19554], bl[19555], bl[19556], bl[19557], bl[19558], bl[19559], bl[19560], bl[19561], bl[19562], bl[19563], bl[19564], bl[19565], bl[19566], bl[19567], bl[19568], bl[19569], bl[19570], bl[19571], bl[19572], bl[19573], bl[19574], bl[19575], bl[19576], bl[19577], bl[19578], bl[19579], bl[19580], bl[19581], bl[19582], bl[19583], bl[19584], bl[19585], bl[19586], bl[19587], bl[19588], bl[19589], bl[19590], bl[19591], bl[19592], bl[19593], bl[19594], bl[19595], bl[19596], bl[19597], bl[19598], bl[19599], bl[19600], bl[19601], bl[19602], bl[19603], bl[19604], bl[19605], bl[19606], bl[19607], bl[19608], bl[19609], bl[19610], bl[19611], bl[19612], bl[19613], bl[19614], bl[19615], bl[19616], bl[19617], bl[19618], bl[19619], bl[19620], bl[19621], bl[19622], bl[19623], bl[19624], bl[19625], bl[19626], bl[19627], bl[19628], bl[19629], bl[19630], bl[19631], bl[19632], bl[19633], bl[19634], bl[19635], bl[19636], bl[19637], bl[19638], bl[19639], bl[19640], bl[19641], bl[19642], bl[19643], bl[19644], bl[19645], bl[19646], bl[19647], bl[19648], bl[19649], bl[19650], bl[19651], bl[19652], bl[19653], bl[19654], bl[19655], bl[19656], bl[19657], bl[19658], bl[19659], bl[19660], bl[19661], bl[19662], bl[19663], bl[19664], bl[19665], bl[19666], bl[19667], bl[19668], bl[19669], bl[19670], bl[19671], bl[19672], bl[19673], bl[19674], bl[19675], bl[19676], bl[19677], bl[19678], bl[19679], bl[19680], bl[19681], bl[19682], bl[19683], bl[19684], bl[19685], bl[19686], bl[19687], bl[19688], bl[19689], bl[19690], bl[19691], bl[19692], bl[19693], bl[19694], bl[19695], bl[19696], bl[19697], bl[19698], bl[19699], bl[19700], bl[19701], bl[19702], bl[19703], bl[19704], bl[19705], bl[19706], bl[19707], bl[19708], bl[19709], bl[19710], bl[19711], bl[19712], bl[19713], bl[19714], bl[19715], bl[19716], bl[19717], bl[19718], bl[19719], bl[19720], bl[19721], bl[19722], bl[19723], bl[19724], bl[19725], bl[19726], bl[19727], bl[19728], bl[19729], bl[19730], bl[19731], bl[19732], bl[19733], bl[19734], bl[19735], bl[19736], bl[19737], bl[19738], bl[19739], bl[19740], bl[19741], bl[19742], bl[19743], bl[19744], bl[19745], bl[19746], bl[19747], bl[19748], bl[19749], bl[19750], bl[19751], bl[19752], bl[19753], bl[19754], bl[19755], bl[19756], bl[19757], bl[19758], bl[19759], bl[19760], bl[19761], bl[19762], bl[19763], bl[19764], bl[19765], bl[19766], bl[19767], bl[19768], bl[19769], bl[19770], bl[19771], bl[19772], bl[19773], bl[19774], bl[19775], bl[19776], bl[19777], bl[19778], bl[19779], bl[19780], bl[19781], bl[19782], bl[19783], bl[19784], bl[19785], bl[19786], bl[19787], bl[19788], bl[19789], bl[19790], bl[19791], bl[19792], bl[19793], bl[19794], bl[19795], bl[19796], bl[19797], bl[19798], bl[19799], bl[19800], bl[19801], bl[19802], bl[19803], bl[19804], bl[19805], bl[19806], bl[19807], bl[19808], bl[19809], bl[19810], bl[19811], bl[19812], bl[19813], bl[19814], bl[19815], bl[19816], bl[19817], bl[19818], bl[19819], bl[19820], bl[19821], bl[19822], bl[19823], bl[19824], bl[19825], bl[19826], bl[19827], bl[19828], bl[19829], bl[19830], bl[19831], bl[19832], bl[19833], bl[19834], bl[19835], bl[19836], bl[19837], bl[19838], bl[19839], bl[19840], bl[19841], bl[19842], bl[19843], bl[19844], bl[19845], bl[19846], bl[19847], bl[19848], bl[19849], bl[19850], bl[19851], bl[19852], bl[19853], bl[19854], bl[19855], bl[19856], bl[19857], bl[19858], bl[19859], bl[19860], bl[19861], bl[19862], bl[19863], bl[19864], bl[19865], bl[19866], bl[19867], bl[19868], bl[19869], bl[19870], bl[19871], bl[19872], bl[19873], bl[19874], bl[19875], bl[19876], bl[19877], bl[19878], bl[19879], bl[19880], bl[19881], bl[19882], bl[19883], bl[19884], bl[19885], bl[19886], bl[19887], bl[19888], bl[19889], bl[19890], bl[19891], bl[19892], bl[19893], bl[19894], bl[19895], bl[19896], bl[19897], bl[19898], bl[19899], bl[19900], bl[19901], bl[19902], bl[19903], bl[19904], bl[19905], bl[19906], bl[19907], bl[19908], bl[19909], bl[19910], bl[19911], bl[19912], bl[19913], bl[19914], bl[19915], bl[19916], bl[19917], bl[19918], bl[19919], bl[19920], bl[19921], bl[19922], bl[19923], bl[19924], bl[19925], bl[19926], bl[19927], bl[19928], bl[19929], bl[19930], bl[19931], bl[19932], bl[19933], bl[19934], bl[19935], bl[19936], bl[19937], bl[19938], bl[19939], bl[19940], bl[19941], bl[19942], bl[19943], bl[19944], bl[19945], bl[19946], bl[19947], bl[19948], bl[19949], bl[19950], bl[19951], bl[19952], bl[19953], bl[19954], bl[19955], bl[19956], bl[19957], bl[19958], bl[19959], bl[19960], bl[19961], bl[19962], bl[19963], bl[19964], bl[19965], bl[19966], bl[19967], bl[19968], bl[19969], bl[19970], bl[19971], bl[19972], bl[19973], bl[19974], bl[19975], bl[19976], bl[19977], bl[19978], bl[19979], bl[19980], bl[19981], bl[19982], bl[19983], bl[19984], bl[19985], bl[19986], bl[19987], bl[19988], bl[19989], bl[19990], bl[19991], bl[19992], bl[19993], bl[19994], bl[19995], bl[19996], bl[19997], bl[19998], bl[19999], bl[20000], bl[20001], bl[20002], bl[20003], bl[20004], bl[20005], bl[20006], bl[20007], bl[20008], bl[20009], bl[20010], bl[20011], bl[20012], bl[20013], bl[20014], bl[20015], bl[20016], bl[20017], bl[20018], bl[20019], bl[20020], bl[20021], bl[20022], bl[20023], bl[20024], bl[20025], bl[20026], bl[20027], bl[20028], bl[20029], bl[20030], bl[20031], bl[20032], bl[20033], bl[20034], bl[20035], bl[20036], bl[20037], bl[20038], bl[20039], bl[20040], bl[20041], bl[20042], bl[20043], bl[20044], bl[20045], bl[20046], bl[20047], bl[20048], bl[20049], bl[20050], bl[20051], bl[20052], bl[20053], bl[20054], bl[20055], bl[20056], bl[20057], bl[20058], bl[20059], bl[20060], bl[20061], bl[20062], bl[20063], bl[20064], bl[20065], bl[20066], bl[20067], bl[20068], bl[20069], bl[20070], bl[20071], bl[20072], bl[20073], bl[20074], bl[20075], bl[20076], bl[20077], bl[20078], bl[20079], bl[20080], bl[20081], bl[20082], bl[20083], bl[20084], bl[20085], bl[20086], bl[20087], bl[20088], bl[20089], bl[20090], bl[20091], bl[20092], bl[20093], bl[20094], bl[20095], bl[20096], bl[20097], bl[20098], bl[20099], bl[20100], bl[20101], bl[20102], bl[20103], bl[20104], bl[20105], bl[20106], bl[20107], bl[20108], bl[20109], bl[20110], bl[20111], bl[20112], bl[20113], bl[20114], bl[20115], bl[20116], bl[20117], bl[20118], bl[20119], bl[20120], bl[20121], bl[20122], bl[20123], bl[20124], bl[20125], bl[20126], bl[20127], bl[20128], bl[20129], bl[20130], bl[20131], bl[20132], bl[20133], bl[20134], bl[20135], bl[20136], bl[20137], bl[20138], bl[20139], bl[20140], bl[20141], bl[20142], bl[20143], bl[20144], bl[20145], bl[20146], bl[20147], bl[20148], bl[20149], bl[20150], bl[20151], bl[20152], bl[20153], bl[20154], bl[20155], bl[20156], bl[20157], bl[20158], bl[20159], bl[20160], bl[20161], bl[20162], bl[20163], bl[20164], bl[20165], bl[20166], bl[20167], bl[20168], bl[20169], bl[20170], bl[20171], bl[20172], bl[20173], bl[20174], bl[20175], bl[20176], bl[20177], bl[20178], bl[20179], bl[20180], bl[20181], bl[20182], bl[20183], bl[20184], bl[20185], bl[20186], bl[20187], bl[20188], bl[20189], bl[20190], bl[20191], bl[20192], bl[20193], bl[20194], bl[20195], bl[20196], bl[20197], bl[20198], bl[20199], bl[20200], bl[20201], bl[20202], bl[20203], bl[20204], bl[20205], bl[20206], bl[20207], bl[20208], bl[20209], bl[20210], bl[20211], bl[20212], bl[20213], bl[20214], bl[20215], bl[20216], bl[20217], bl[20218], bl[20219], bl[20220], bl[20221], bl[20222], bl[20223], bl[20224], bl[20225], bl[20226], bl[20227], bl[20228], bl[20229], bl[20230], bl[20231], bl[20232], bl[20233], bl[20234], bl[20235], bl[20236], bl[20237], bl[20238], bl[20239], bl[20240], bl[20241], bl[20242], bl[20243], bl[20244], bl[20245], bl[20246], bl[20247], bl[536], bl[537], bl[538], bl[539], bl[540], bl[541], bl[542], bl[543], bl[464], bl[465], bl[466], bl[467], bl[468], bl[469], bl[470], bl[471], bl[472], bl[473], bl[474], bl[475], bl[476], bl[477], bl[478], bl[479], bl[480], bl[481], bl[482], bl[483], bl[484], bl[485], bl[486], bl[487], bl[488], bl[489], bl[490], bl[491], bl[492], bl[493], bl[494], bl[495], bl[496], bl[497], bl[498], bl[499], bl[500], bl[501], bl[502], bl[503], bl[504], bl[505], bl[506], bl[507], bl[508], bl[509], bl[510], bl[511], bl[512], bl[513], bl[514], bl[515], bl[516], bl[517], bl[518], bl[519], bl[520], bl[521], bl[522], bl[523], bl[524], bl[525], bl[526], bl[527], bl[528], bl[529], bl[530], bl[531], bl[532], bl[533], bl[534], bl[535], bl[19148], bl[19149], bl[19150], bl[19151], bl[19152], bl[19153], bl[19154], bl[19155], bl[19156], bl[19157], bl[19158], bl[19159], bl[19160], bl[19161], bl[19162], bl[19163], bl[19164], bl[19165], bl[19166], bl[19167], bl[19168], bl[19169], bl[19170], bl[19171], bl[19172], bl[19173], bl[19174], bl[19175], bl[19176], bl[19177], bl[19178], bl[19179], bl[19180], bl[19181], bl[19182], bl[19183], bl[19184], bl[19185], bl[19186], bl[19187], bl[19188], bl[19189], bl[19190], bl[19191], bl[19192], bl[19193], bl[19194], bl[19195], bl[19196], bl[19197], bl[19198], bl[19199], bl[19200], bl[19201], bl[19202], bl[19203], bl[19204], bl[19205], bl[19206], bl[19207], bl[19208], bl[19209], bl[19210], bl[19211], bl[19212], bl[19213], bl[19214], bl[19215], bl[19216], bl[19217], bl[19218], bl[19219], bl[19220], bl[19221], bl[19222], bl[19223], bl[19224], bl[19225], bl[19226], bl[19227], bl[384], bl[385], bl[386], bl[387], bl[388], bl[389], bl[390], bl[391], bl[392], bl[393], bl[394], bl[395], bl[396], bl[397], bl[398], bl[399], bl[400], bl[401], bl[402], bl[403], bl[404], bl[405], bl[406], bl[407], bl[408], bl[409], bl[410], bl[411], bl[412], bl[413], bl[414], bl[415], bl[416], bl[417], bl[418], bl[419], bl[420], bl[421], bl[422], bl[423], bl[424], bl[425], bl[426], bl[427], bl[428], bl[429], bl[430], bl[431], bl[432], bl[433], bl[434], bl[435], bl[436], bl[437], bl[438], bl[439], bl[440], bl[441], bl[442], bl[443], bl[444], bl[445], bl[446], bl[447], bl[448], bl[449], bl[450], bl[451], bl[452], bl[453], bl[454], bl[455], bl[456], bl[457], bl[458], bl[459], bl[460], bl[461], bl[462], bl[463]}),
        .wl({wl[19228], wl[19229], wl[19230], wl[19231], wl[19232], wl[19233], wl[19234], wl[19235], wl[19236], wl[19237], wl[19238], wl[19239], wl[19240], wl[19241], wl[19242], wl[19243], wl[19244], wl[19245], wl[19246], wl[19247], wl[19248], wl[19249], wl[19250], wl[19251], wl[19252], wl[19253], wl[19254], wl[19255], wl[19256], wl[19257], wl[19258], wl[19259], wl[19260], wl[19261], wl[19262], wl[19263], wl[19264], wl[19265], wl[19266], wl[19267], wl[19268], wl[19269], wl[19270], wl[19271], wl[19272], wl[19273], wl[19274], wl[19275], wl[19276], wl[19277], wl[19278], wl[19279], wl[19280], wl[19281], wl[19282], wl[19283], wl[19284], wl[19285], wl[19286], wl[19287], wl[19288], wl[19289], wl[19290], wl[19291], wl[19292], wl[19293], wl[19294], wl[19295], wl[19296], wl[19297], wl[19298], wl[19299], wl[19300], wl[19301], wl[19302], wl[19303], wl[19304], wl[19305], wl[19306], wl[19307], wl[19308], wl[19309], wl[19310], wl[19311], wl[19312], wl[19313], wl[19314], wl[19315], wl[19316], wl[19317], wl[19318], wl[19319], wl[19320], wl[19321], wl[19322], wl[19323], wl[19324], wl[19325], wl[19326], wl[19327], wl[19328], wl[19329], wl[19330], wl[19331], wl[19332], wl[19333], wl[19334], wl[19335], wl[19336], wl[19337], wl[19338], wl[19339], wl[19340], wl[19341], wl[19342], wl[19343], wl[19344], wl[19345], wl[19346], wl[19347], wl[19348], wl[19349], wl[19350], wl[19351], wl[19352], wl[19353], wl[19354], wl[19355], wl[19356], wl[19357], wl[19358], wl[19359], wl[19360], wl[19361], wl[19362], wl[19363], wl[19364], wl[19365], wl[19366], wl[19367], wl[19368], wl[19369], wl[19370], wl[19371], wl[19372], wl[19373], wl[19374], wl[19375], wl[19376], wl[19377], wl[19378], wl[19379], wl[19380], wl[19381], wl[19382], wl[19383], wl[19384], wl[19385], wl[19386], wl[19387], wl[19388], wl[19389], wl[19390], wl[19391], wl[19392], wl[19393], wl[19394], wl[19395], wl[19396], wl[19397], wl[19398], wl[19399], wl[19400], wl[19401], wl[19402], wl[19403], wl[19404], wl[19405], wl[19406], wl[19407], wl[19408], wl[19409], wl[19410], wl[19411], wl[19412], wl[19413], wl[19414], wl[19415], wl[19416], wl[19417], wl[19418], wl[19419], wl[19420], wl[19421], wl[19422], wl[19423], wl[19424], wl[19425], wl[19426], wl[19427], wl[19428], wl[19429], wl[19430], wl[19431], wl[19432], wl[19433], wl[19434], wl[19435], wl[19436], wl[19437], wl[19438], wl[19439], wl[19440], wl[19441], wl[19442], wl[19443], wl[19444], wl[19445], wl[19446], wl[19447], wl[19448], wl[19449], wl[19450], wl[19451], wl[19452], wl[19453], wl[19454], wl[19455], wl[19456], wl[19457], wl[19458], wl[19459], wl[19460], wl[19461], wl[19462], wl[19463], wl[19464], wl[19465], wl[19466], wl[19467], wl[19468], wl[19469], wl[19470], wl[19471], wl[19472], wl[19473], wl[19474], wl[19475], wl[19476], wl[19477], wl[19478], wl[19479], wl[19480], wl[19481], wl[19482], wl[19483], wl[19484], wl[19485], wl[19486], wl[19487], wl[19488], wl[19489], wl[19490], wl[19491], wl[19492], wl[19493], wl[19494], wl[19495], wl[19496], wl[19497], wl[19498], wl[19499], wl[19500], wl[19501], wl[19502], wl[19503], wl[19504], wl[19505], wl[19506], wl[19507], wl[19508], wl[19509], wl[19510], wl[19511], wl[19512], wl[19513], wl[19514], wl[19515], wl[19516], wl[19517], wl[19518], wl[19519], wl[19520], wl[19521], wl[19522], wl[19523], wl[19524], wl[19525], wl[19526], wl[19527], wl[19528], wl[19529], wl[19530], wl[19531], wl[19532], wl[19533], wl[19534], wl[19535], wl[19536], wl[19537], wl[19538], wl[19539], wl[19540], wl[19541], wl[19542], wl[19543], wl[19544], wl[19545], wl[19546], wl[19547], wl[19548], wl[19549], wl[19550], wl[19551], wl[19552], wl[19553], wl[19554], wl[19555], wl[19556], wl[19557], wl[19558], wl[19559], wl[19560], wl[19561], wl[19562], wl[19563], wl[19564], wl[19565], wl[19566], wl[19567], wl[19568], wl[19569], wl[19570], wl[19571], wl[19572], wl[19573], wl[19574], wl[19575], wl[19576], wl[19577], wl[19578], wl[19579], wl[19580], wl[19581], wl[19582], wl[19583], wl[19584], wl[19585], wl[19586], wl[19587], wl[19588], wl[19589], wl[19590], wl[19591], wl[19592], wl[19593], wl[19594], wl[19595], wl[19596], wl[19597], wl[19598], wl[19599], wl[19600], wl[19601], wl[19602], wl[19603], wl[19604], wl[19605], wl[19606], wl[19607], wl[19608], wl[19609], wl[19610], wl[19611], wl[19612], wl[19613], wl[19614], wl[19615], wl[19616], wl[19617], wl[19618], wl[19619], wl[19620], wl[19621], wl[19622], wl[19623], wl[19624], wl[19625], wl[19626], wl[19627], wl[19628], wl[19629], wl[19630], wl[19631], wl[19632], wl[19633], wl[19634], wl[19635], wl[19636], wl[19637], wl[19638], wl[19639], wl[19640], wl[19641], wl[19642], wl[19643], wl[19644], wl[19645], wl[19646], wl[19647], wl[19648], wl[19649], wl[19650], wl[19651], wl[19652], wl[19653], wl[19654], wl[19655], wl[19656], wl[19657], wl[19658], wl[19659], wl[19660], wl[19661], wl[19662], wl[19663], wl[19664], wl[19665], wl[19666], wl[19667], wl[19668], wl[19669], wl[19670], wl[19671], wl[19672], wl[19673], wl[19674], wl[19675], wl[19676], wl[19677], wl[19678], wl[19679], wl[19680], wl[19681], wl[19682], wl[19683], wl[19684], wl[19685], wl[19686], wl[19687], wl[19688], wl[19689], wl[19690], wl[19691], wl[19692], wl[19693], wl[19694], wl[19695], wl[19696], wl[19697], wl[19698], wl[19699], wl[19700], wl[19701], wl[19702], wl[19703], wl[19704], wl[19705], wl[19706], wl[19707], wl[19708], wl[19709], wl[19710], wl[19711], wl[19712], wl[19713], wl[19714], wl[19715], wl[19716], wl[19717], wl[19718], wl[19719], wl[19720], wl[19721], wl[19722], wl[19723], wl[19724], wl[19725], wl[19726], wl[19727], wl[19728], wl[19729], wl[19730], wl[19731], wl[19732], wl[19733], wl[19734], wl[19735], wl[19736], wl[19737], wl[19738], wl[19739], wl[19740], wl[19741], wl[19742], wl[19743], wl[19744], wl[19745], wl[19746], wl[19747], wl[19748], wl[19749], wl[19750], wl[19751], wl[19752], wl[19753], wl[19754], wl[19755], wl[19756], wl[19757], wl[19758], wl[19759], wl[19760], wl[19761], wl[19762], wl[19763], wl[19764], wl[19765], wl[19766], wl[19767], wl[19768], wl[19769], wl[19770], wl[19771], wl[19772], wl[19773], wl[19774], wl[19775], wl[19776], wl[19777], wl[19778], wl[19779], wl[19780], wl[19781], wl[19782], wl[19783], wl[19784], wl[19785], wl[19786], wl[19787], wl[19788], wl[19789], wl[19790], wl[19791], wl[19792], wl[19793], wl[19794], wl[19795], wl[19796], wl[19797], wl[19798], wl[19799], wl[19800], wl[19801], wl[19802], wl[19803], wl[19804], wl[19805], wl[19806], wl[19807], wl[19808], wl[19809], wl[19810], wl[19811], wl[19812], wl[19813], wl[19814], wl[19815], wl[19816], wl[19817], wl[19818], wl[19819], wl[19820], wl[19821], wl[19822], wl[19823], wl[19824], wl[19825], wl[19826], wl[19827], wl[19828], wl[19829], wl[19830], wl[19831], wl[19832], wl[19833], wl[19834], wl[19835], wl[19836], wl[19837], wl[19838], wl[19839], wl[19840], wl[19841], wl[19842], wl[19843], wl[19844], wl[19845], wl[19846], wl[19847], wl[19848], wl[19849], wl[19850], wl[19851], wl[19852], wl[19853], wl[19854], wl[19855], wl[19856], wl[19857], wl[19858], wl[19859], wl[19860], wl[19861], wl[19862], wl[19863], wl[19864], wl[19865], wl[19866], wl[19867], wl[19868], wl[19869], wl[19870], wl[19871], wl[19872], wl[19873], wl[19874], wl[19875], wl[19876], wl[19877], wl[19878], wl[19879], wl[19880], wl[19881], wl[19882], wl[19883], wl[19884], wl[19885], wl[19886], wl[19887], wl[19888], wl[19889], wl[19890], wl[19891], wl[19892], wl[19893], wl[19894], wl[19895], wl[19896], wl[19897], wl[19898], wl[19899], wl[19900], wl[19901], wl[19902], wl[19903], wl[19904], wl[19905], wl[19906], wl[19907], wl[19908], wl[19909], wl[19910], wl[19911], wl[19912], wl[19913], wl[19914], wl[19915], wl[19916], wl[19917], wl[19918], wl[19919], wl[19920], wl[19921], wl[19922], wl[19923], wl[19924], wl[19925], wl[19926], wl[19927], wl[19928], wl[19929], wl[19930], wl[19931], wl[19932], wl[19933], wl[19934], wl[19935], wl[19936], wl[19937], wl[19938], wl[19939], wl[19940], wl[19941], wl[19942], wl[19943], wl[19944], wl[19945], wl[19946], wl[19947], wl[19948], wl[19949], wl[19950], wl[19951], wl[19952], wl[19953], wl[19954], wl[19955], wl[19956], wl[19957], wl[19958], wl[19959], wl[19960], wl[19961], wl[19962], wl[19963], wl[19964], wl[19965], wl[19966], wl[19967], wl[19968], wl[19969], wl[19970], wl[19971], wl[19972], wl[19973], wl[19974], wl[19975], wl[19976], wl[19977], wl[19978], wl[19979], wl[19980], wl[19981], wl[19982], wl[19983], wl[19984], wl[19985], wl[19986], wl[19987], wl[19988], wl[19989], wl[19990], wl[19991], wl[19992], wl[19993], wl[19994], wl[19995], wl[19996], wl[19997], wl[19998], wl[19999], wl[20000], wl[20001], wl[20002], wl[20003], wl[20004], wl[20005], wl[20006], wl[20007], wl[20008], wl[20009], wl[20010], wl[20011], wl[20012], wl[20013], wl[20014], wl[20015], wl[20016], wl[20017], wl[20018], wl[20019], wl[20020], wl[20021], wl[20022], wl[20023], wl[20024], wl[20025], wl[20026], wl[20027], wl[20028], wl[20029], wl[20030], wl[20031], wl[20032], wl[20033], wl[20034], wl[20035], wl[20036], wl[20037], wl[20038], wl[20039], wl[20040], wl[20041], wl[20042], wl[20043], wl[20044], wl[20045], wl[20046], wl[20047], wl[20048], wl[20049], wl[20050], wl[20051], wl[20052], wl[20053], wl[20054], wl[20055], wl[20056], wl[20057], wl[20058], wl[20059], wl[20060], wl[20061], wl[20062], wl[20063], wl[20064], wl[20065], wl[20066], wl[20067], wl[20068], wl[20069], wl[20070], wl[20071], wl[20072], wl[20073], wl[20074], wl[20075], wl[20076], wl[20077], wl[20078], wl[20079], wl[20080], wl[20081], wl[20082], wl[20083], wl[20084], wl[20085], wl[20086], wl[20087], wl[20088], wl[20089], wl[20090], wl[20091], wl[20092], wl[20093], wl[20094], wl[20095], wl[20096], wl[20097], wl[20098], wl[20099], wl[20100], wl[20101], wl[20102], wl[20103], wl[20104], wl[20105], wl[20106], wl[20107], wl[20108], wl[20109], wl[20110], wl[20111], wl[20112], wl[20113], wl[20114], wl[20115], wl[20116], wl[20117], wl[20118], wl[20119], wl[20120], wl[20121], wl[20122], wl[20123], wl[20124], wl[20125], wl[20126], wl[20127], wl[20128], wl[20129], wl[20130], wl[20131], wl[20132], wl[20133], wl[20134], wl[20135], wl[20136], wl[20137], wl[20138], wl[20139], wl[20140], wl[20141], wl[20142], wl[20143], wl[20144], wl[20145], wl[20146], wl[20147], wl[20148], wl[20149], wl[20150], wl[20151], wl[20152], wl[20153], wl[20154], wl[20155], wl[20156], wl[20157], wl[20158], wl[20159], wl[20160], wl[20161], wl[20162], wl[20163], wl[20164], wl[20165], wl[20166], wl[20167], wl[20168], wl[20169], wl[20170], wl[20171], wl[20172], wl[20173], wl[20174], wl[20175], wl[20176], wl[20177], wl[20178], wl[20179], wl[20180], wl[20181], wl[20182], wl[20183], wl[20184], wl[20185], wl[20186], wl[20187], wl[20188], wl[20189], wl[20190], wl[20191], wl[20192], wl[20193], wl[20194], wl[20195], wl[20196], wl[20197], wl[20198], wl[20199], wl[20200], wl[20201], wl[20202], wl[20203], wl[20204], wl[20205], wl[20206], wl[20207], wl[20208], wl[20209], wl[20210], wl[20211], wl[20212], wl[20213], wl[20214], wl[20215], wl[20216], wl[20217], wl[20218], wl[20219], wl[20220], wl[20221], wl[20222], wl[20223], wl[20224], wl[20225], wl[20226], wl[20227], wl[20228], wl[20229], wl[20230], wl[20231], wl[20232], wl[20233], wl[20234], wl[20235], wl[20236], wl[20237], wl[20238], wl[20239], wl[20240], wl[20241], wl[20242], wl[20243], wl[20244], wl[20245], wl[20246], wl[20247], wl[536], wl[537], wl[538], wl[539], wl[540], wl[541], wl[542], wl[543], wl[464], wl[465], wl[466], wl[467], wl[468], wl[469], wl[470], wl[471], wl[472], wl[473], wl[474], wl[475], wl[476], wl[477], wl[478], wl[479], wl[480], wl[481], wl[482], wl[483], wl[484], wl[485], wl[486], wl[487], wl[488], wl[489], wl[490], wl[491], wl[492], wl[493], wl[494], wl[495], wl[496], wl[497], wl[498], wl[499], wl[500], wl[501], wl[502], wl[503], wl[504], wl[505], wl[506], wl[507], wl[508], wl[509], wl[510], wl[511], wl[512], wl[513], wl[514], wl[515], wl[516], wl[517], wl[518], wl[519], wl[520], wl[521], wl[522], wl[523], wl[524], wl[525], wl[526], wl[527], wl[528], wl[529], wl[530], wl[531], wl[532], wl[533], wl[534], wl[535], wl[19148], wl[19149], wl[19150], wl[19151], wl[19152], wl[19153], wl[19154], wl[19155], wl[19156], wl[19157], wl[19158], wl[19159], wl[19160], wl[19161], wl[19162], wl[19163], wl[19164], wl[19165], wl[19166], wl[19167], wl[19168], wl[19169], wl[19170], wl[19171], wl[19172], wl[19173], wl[19174], wl[19175], wl[19176], wl[19177], wl[19178], wl[19179], wl[19180], wl[19181], wl[19182], wl[19183], wl[19184], wl[19185], wl[19186], wl[19187], wl[19188], wl[19189], wl[19190], wl[19191], wl[19192], wl[19193], wl[19194], wl[19195], wl[19196], wl[19197], wl[19198], wl[19199], wl[19200], wl[19201], wl[19202], wl[19203], wl[19204], wl[19205], wl[19206], wl[19207], wl[19208], wl[19209], wl[19210], wl[19211], wl[19212], wl[19213], wl[19214], wl[19215], wl[19216], wl[19217], wl[19218], wl[19219], wl[19220], wl[19221], wl[19222], wl[19223], wl[19224], wl[19225], wl[19226], wl[19227], wl[384], wl[385], wl[386], wl[387], wl[388], wl[389], wl[390], wl[391], wl[392], wl[393], wl[394], wl[395], wl[396], wl[397], wl[398], wl[399], wl[400], wl[401], wl[402], wl[403], wl[404], wl[405], wl[406], wl[407], wl[408], wl[409], wl[410], wl[411], wl[412], wl[413], wl[414], wl[415], wl[416], wl[417], wl[418], wl[419], wl[420], wl[421], wl[422], wl[423], wl[424], wl[425], wl[426], wl[427], wl[428], wl[429], wl[430], wl[431], wl[432], wl[433], wl[434], wl[435], wl[436], wl[437], wl[438], wl[439], wl[440], wl[441], wl[442], wl[443], wl[444], wl[445], wl[446], wl[447], wl[448], wl[449], wl[450], wl[451], wl[452], wl[453], wl[454], wl[455], wl[456], wl[457], wl[458], wl[459], wl[460], wl[461], wl[462], wl[463]})
    );
    top_tile tile_4__5_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_2__4__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_2__4__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_2__4__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_3__3__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_3__3__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_3__3__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_2__3__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_2__3__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_2__3__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_2__3__grid_top_r_in[1]),
        .grid_left_in(grid_clb_3__4__grid_left_in),
        .grid_bottom_in(grid_clb_3__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[16:23]),
        .io_bottom_in(grid_io_top_3__5__io_bottom_in),
        .chanx_left_in(sb_1__4__1_chanx_right_out),
        .chanx_left_out(cbx_1__4__2_chanx_left_out),
        .chany_bottom_in(sb_1__1__8_chany_top_out),
        .chany_bottom_out(cby_1__1__11_chany_bottom_out),
        .grid_right_out(grid_clb_4__4__grid_left_in),
        .chanx_right_in_0(cbx_1__4__3_chanx_left_out),
        .chanx_right_out_0(sb_1__4__2_chanx_right_out),
        .grid_right_t_inpad(grid_io_top_4__5__io_bottom_in),
        .grid_right_b_in(sb_3__4__grid_right_b_in),
        .grid_bottom_r_in(sb_3__3__grid_top_r_in),
        .grid_bottom_l_in(sb_3__3__grid_top_l_in),
        .grid_left_b_in(sb_2__4__grid_right_b_in),
        .bl({bl[17968], bl[17969], bl[17970], bl[17971], bl[17972], bl[17973], bl[17974], bl[17975], bl[17976], bl[17977], bl[17978], bl[17979], bl[17980], bl[17981], bl[17982], bl[17983], bl[17984], bl[17985], bl[17986], bl[17987], bl[17988], bl[17989], bl[17990], bl[17991], bl[17992], bl[17993], bl[17994], bl[17995], bl[17996], bl[17997], bl[17998], bl[17999], bl[18000], bl[18001], bl[18002], bl[18003], bl[18004], bl[18005], bl[18006], bl[18007], bl[18008], bl[18009], bl[18010], bl[18011], bl[18012], bl[18013], bl[18014], bl[18015], bl[18016], bl[18017], bl[18018], bl[18019], bl[18020], bl[18021], bl[18022], bl[18023], bl[18024], bl[18025], bl[18026], bl[18027], bl[18028], bl[18029], bl[18030], bl[18031], bl[18032], bl[18033], bl[18034], bl[18035], bl[18036], bl[18037], bl[18038], bl[18039], bl[18040], bl[18041], bl[18042], bl[18043], bl[18044], bl[18045], bl[18046], bl[18047], bl[18048], bl[18049], bl[18050], bl[18051], bl[18052], bl[18053], bl[18054], bl[18055], bl[18056], bl[18057], bl[18058], bl[18059], bl[18060], bl[18061], bl[18062], bl[18063], bl[18064], bl[18065], bl[18066], bl[18067], bl[18068], bl[18069], bl[18070], bl[18071], bl[18072], bl[18073], bl[18074], bl[18075], bl[18076], bl[18077], bl[18078], bl[18079], bl[18080], bl[18081], bl[18082], bl[18083], bl[18084], bl[18085], bl[18086], bl[18087], bl[18088], bl[18089], bl[18090], bl[18091], bl[18092], bl[18093], bl[18094], bl[18095], bl[18096], bl[18097], bl[18098], bl[18099], bl[18100], bl[18101], bl[18102], bl[18103], bl[18104], bl[18105], bl[18106], bl[18107], bl[18108], bl[18109], bl[18110], bl[18111], bl[18112], bl[18113], bl[18114], bl[18115], bl[18116], bl[18117], bl[18118], bl[18119], bl[18120], bl[18121], bl[18122], bl[18123], bl[18124], bl[18125], bl[18126], bl[18127], bl[18128], bl[18129], bl[18130], bl[18131], bl[18132], bl[18133], bl[18134], bl[18135], bl[18136], bl[18137], bl[18138], bl[18139], bl[18140], bl[18141], bl[18142], bl[18143], bl[18144], bl[18145], bl[18146], bl[18147], bl[18148], bl[18149], bl[18150], bl[18151], bl[18152], bl[18153], bl[18154], bl[18155], bl[18156], bl[18157], bl[18158], bl[18159], bl[18160], bl[18161], bl[18162], bl[18163], bl[18164], bl[18165], bl[18166], bl[18167], bl[18168], bl[18169], bl[18170], bl[18171], bl[18172], bl[18173], bl[18174], bl[18175], bl[18176], bl[18177], bl[18178], bl[18179], bl[18180], bl[18181], bl[18182], bl[18183], bl[18184], bl[18185], bl[18186], bl[18187], bl[18188], bl[18189], bl[18190], bl[18191], bl[18192], bl[18193], bl[18194], bl[18195], bl[18196], bl[18197], bl[18198], bl[18199], bl[18200], bl[18201], bl[18202], bl[18203], bl[18204], bl[18205], bl[18206], bl[18207], bl[18208], bl[18209], bl[18210], bl[18211], bl[18212], bl[18213], bl[18214], bl[18215], bl[18216], bl[18217], bl[18218], bl[18219], bl[18220], bl[18221], bl[18222], bl[18223], bl[18224], bl[18225], bl[18226], bl[18227], bl[18228], bl[18229], bl[18230], bl[18231], bl[18232], bl[18233], bl[18234], bl[18235], bl[18236], bl[18237], bl[18238], bl[18239], bl[18240], bl[18241], bl[18242], bl[18243], bl[18244], bl[18245], bl[18246], bl[18247], bl[18248], bl[18249], bl[18250], bl[18251], bl[18252], bl[18253], bl[18254], bl[18255], bl[18256], bl[18257], bl[18258], bl[18259], bl[18260], bl[18261], bl[18262], bl[18263], bl[18264], bl[18265], bl[18266], bl[18267], bl[18268], bl[18269], bl[18270], bl[18271], bl[18272], bl[18273], bl[18274], bl[18275], bl[18276], bl[18277], bl[18278], bl[18279], bl[18280], bl[18281], bl[18282], bl[18283], bl[18284], bl[18285], bl[18286], bl[18287], bl[18288], bl[18289], bl[18290], bl[18291], bl[18292], bl[18293], bl[18294], bl[18295], bl[18296], bl[18297], bl[18298], bl[18299], bl[18300], bl[18301], bl[18302], bl[18303], bl[18304], bl[18305], bl[18306], bl[18307], bl[18308], bl[18309], bl[18310], bl[18311], bl[18312], bl[18313], bl[18314], bl[18315], bl[18316], bl[18317], bl[18318], bl[18319], bl[18320], bl[18321], bl[18322], bl[18323], bl[18324], bl[18325], bl[18326], bl[18327], bl[18328], bl[18329], bl[18330], bl[18331], bl[18332], bl[18333], bl[18334], bl[18335], bl[18336], bl[18337], bl[18338], bl[18339], bl[18340], bl[18341], bl[18342], bl[18343], bl[18344], bl[18345], bl[18346], bl[18347], bl[18348], bl[18349], bl[18350], bl[18351], bl[18352], bl[18353], bl[18354], bl[18355], bl[18356], bl[18357], bl[18358], bl[18359], bl[18360], bl[18361], bl[18362], bl[18363], bl[18364], bl[18365], bl[18366], bl[18367], bl[18368], bl[18369], bl[18370], bl[18371], bl[18372], bl[18373], bl[18374], bl[18375], bl[18376], bl[18377], bl[18378], bl[18379], bl[18380], bl[18381], bl[18382], bl[18383], bl[18384], bl[18385], bl[18386], bl[18387], bl[18388], bl[18389], bl[18390], bl[18391], bl[18392], bl[18393], bl[18394], bl[18395], bl[18396], bl[18397], bl[18398], bl[18399], bl[18400], bl[18401], bl[18402], bl[18403], bl[18404], bl[18405], bl[18406], bl[18407], bl[18408], bl[18409], bl[18410], bl[18411], bl[18412], bl[18413], bl[18414], bl[18415], bl[18416], bl[18417], bl[18418], bl[18419], bl[18420], bl[18421], bl[18422], bl[18423], bl[18424], bl[18425], bl[18426], bl[18427], bl[18428], bl[18429], bl[18430], bl[18431], bl[18432], bl[18433], bl[18434], bl[18435], bl[18436], bl[18437], bl[18438], bl[18439], bl[18440], bl[18441], bl[18442], bl[18443], bl[18444], bl[18445], bl[18446], bl[18447], bl[18448], bl[18449], bl[18450], bl[18451], bl[18452], bl[18453], bl[18454], bl[18455], bl[18456], bl[18457], bl[18458], bl[18459], bl[18460], bl[18461], bl[18462], bl[18463], bl[18464], bl[18465], bl[18466], bl[18467], bl[18468], bl[18469], bl[18470], bl[18471], bl[18472], bl[18473], bl[18474], bl[18475], bl[18476], bl[18477], bl[18478], bl[18479], bl[18480], bl[18481], bl[18482], bl[18483], bl[18484], bl[18485], bl[18486], bl[18487], bl[18488], bl[18489], bl[18490], bl[18491], bl[18492], bl[18493], bl[18494], bl[18495], bl[18496], bl[18497], bl[18498], bl[18499], bl[18500], bl[18501], bl[18502], bl[18503], bl[18504], bl[18505], bl[18506], bl[18507], bl[18508], bl[18509], bl[18510], bl[18511], bl[18512], bl[18513], bl[18514], bl[18515], bl[18516], bl[18517], bl[18518], bl[18519], bl[18520], bl[18521], bl[18522], bl[18523], bl[18524], bl[18525], bl[18526], bl[18527], bl[18528], bl[18529], bl[18530], bl[18531], bl[18532], bl[18533], bl[18534], bl[18535], bl[18536], bl[18537], bl[18538], bl[18539], bl[18540], bl[18541], bl[18542], bl[18543], bl[18544], bl[18545], bl[18546], bl[18547], bl[18548], bl[18549], bl[18550], bl[18551], bl[18552], bl[18553], bl[18554], bl[18555], bl[18556], bl[18557], bl[18558], bl[18559], bl[18560], bl[18561], bl[18562], bl[18563], bl[18564], bl[18565], bl[18566], bl[18567], bl[18568], bl[18569], bl[18570], bl[18571], bl[18572], bl[18573], bl[18574], bl[18575], bl[18576], bl[18577], bl[18578], bl[18579], bl[18580], bl[18581], bl[18582], bl[18583], bl[18584], bl[18585], bl[18586], bl[18587], bl[18588], bl[18589], bl[18590], bl[18591], bl[18592], bl[18593], bl[18594], bl[18595], bl[18596], bl[18597], bl[18598], bl[18599], bl[18600], bl[18601], bl[18602], bl[18603], bl[18604], bl[18605], bl[18606], bl[18607], bl[18608], bl[18609], bl[18610], bl[18611], bl[18612], bl[18613], bl[18614], bl[18615], bl[18616], bl[18617], bl[18618], bl[18619], bl[18620], bl[18621], bl[18622], bl[18623], bl[18624], bl[18625], bl[18626], bl[18627], bl[18628], bl[18629], bl[18630], bl[18631], bl[18632], bl[18633], bl[18634], bl[18635], bl[18636], bl[18637], bl[18638], bl[18639], bl[18640], bl[18641], bl[18642], bl[18643], bl[18644], bl[18645], bl[18646], bl[18647], bl[18648], bl[18649], bl[18650], bl[18651], bl[18652], bl[18653], bl[18654], bl[18655], bl[18656], bl[18657], bl[18658], bl[18659], bl[18660], bl[18661], bl[18662], bl[18663], bl[18664], bl[18665], bl[18666], bl[18667], bl[18668], bl[18669], bl[18670], bl[18671], bl[18672], bl[18673], bl[18674], bl[18675], bl[18676], bl[18677], bl[18678], bl[18679], bl[18680], bl[18681], bl[18682], bl[18683], bl[18684], bl[18685], bl[18686], bl[18687], bl[18688], bl[18689], bl[18690], bl[18691], bl[18692], bl[18693], bl[18694], bl[18695], bl[18696], bl[18697], bl[18698], bl[18699], bl[18700], bl[18701], bl[18702], bl[18703], bl[18704], bl[18705], bl[18706], bl[18707], bl[18708], bl[18709], bl[18710], bl[18711], bl[18712], bl[18713], bl[18714], bl[18715], bl[18716], bl[18717], bl[18718], bl[18719], bl[18720], bl[18721], bl[18722], bl[18723], bl[18724], bl[18725], bl[18726], bl[18727], bl[18728], bl[18729], bl[18730], bl[18731], bl[18732], bl[18733], bl[18734], bl[18735], bl[18736], bl[18737], bl[18738], bl[18739], bl[18740], bl[18741], bl[18742], bl[18743], bl[18744], bl[18745], bl[18746], bl[18747], bl[18748], bl[18749], bl[18750], bl[18751], bl[18752], bl[18753], bl[18754], bl[18755], bl[18756], bl[18757], bl[18758], bl[18759], bl[18760], bl[18761], bl[18762], bl[18763], bl[18764], bl[18765], bl[18766], bl[18767], bl[18768], bl[18769], bl[18770], bl[18771], bl[18772], bl[18773], bl[18774], bl[18775], bl[18776], bl[18777], bl[18778], bl[18779], bl[18780], bl[18781], bl[18782], bl[18783], bl[18784], bl[18785], bl[18786], bl[18787], bl[18788], bl[18789], bl[18790], bl[18791], bl[18792], bl[18793], bl[18794], bl[18795], bl[18796], bl[18797], bl[18798], bl[18799], bl[18800], bl[18801], bl[18802], bl[18803], bl[18804], bl[18805], bl[18806], bl[18807], bl[18808], bl[18809], bl[18810], bl[18811], bl[18812], bl[18813], bl[18814], bl[18815], bl[18816], bl[18817], bl[18818], bl[18819], bl[18820], bl[18821], bl[18822], bl[18823], bl[18824], bl[18825], bl[18826], bl[18827], bl[18828], bl[18829], bl[18830], bl[18831], bl[18832], bl[18833], bl[18834], bl[18835], bl[18836], bl[18837], bl[18838], bl[18839], bl[18840], bl[18841], bl[18842], bl[18843], bl[18844], bl[18845], bl[18846], bl[18847], bl[18848], bl[18849], bl[18850], bl[18851], bl[18852], bl[18853], bl[18854], bl[18855], bl[18856], bl[18857], bl[18858], bl[18859], bl[18860], bl[18861], bl[18862], bl[18863], bl[18864], bl[18865], bl[18866], bl[18867], bl[18868], bl[18869], bl[18870], bl[18871], bl[18872], bl[18873], bl[18874], bl[18875], bl[18876], bl[18877], bl[18878], bl[18879], bl[18880], bl[18881], bl[18882], bl[18883], bl[18884], bl[18885], bl[18886], bl[18887], bl[18888], bl[18889], bl[18890], bl[18891], bl[18892], bl[18893], bl[18894], bl[18895], bl[18896], bl[18897], bl[18898], bl[18899], bl[18900], bl[18901], bl[18902], bl[18903], bl[18904], bl[18905], bl[18906], bl[18907], bl[18908], bl[18909], bl[18910], bl[18911], bl[18912], bl[18913], bl[18914], bl[18915], bl[18916], bl[18917], bl[18918], bl[18919], bl[18920], bl[18921], bl[18922], bl[18923], bl[18924], bl[18925], bl[18926], bl[18927], bl[18928], bl[18929], bl[18930], bl[18931], bl[18932], bl[18933], bl[18934], bl[18935], bl[18936], bl[18937], bl[18938], bl[18939], bl[18940], bl[18941], bl[18942], bl[18943], bl[18944], bl[18945], bl[18946], bl[18947], bl[18948], bl[18949], bl[18950], bl[18951], bl[18952], bl[18953], bl[18954], bl[18955], bl[18956], bl[18957], bl[18958], bl[18959], bl[18960], bl[18961], bl[18962], bl[18963], bl[18964], bl[18965], bl[18966], bl[18967], bl[18968], bl[18969], bl[18970], bl[18971], bl[18972], bl[18973], bl[18974], bl[18975], bl[18976], bl[18977], bl[18978], bl[18979], bl[18980], bl[18981], bl[18982], bl[18983], bl[18984], bl[18985], bl[18986], bl[18987], bl[376], bl[377], bl[378], bl[379], bl[380], bl[381], bl[382], bl[383], bl[304], bl[305], bl[306], bl[307], bl[308], bl[309], bl[310], bl[311], bl[312], bl[313], bl[314], bl[315], bl[316], bl[317], bl[318], bl[319], bl[320], bl[321], bl[322], bl[323], bl[324], bl[325], bl[326], bl[327], bl[328], bl[329], bl[330], bl[331], bl[332], bl[333], bl[334], bl[335], bl[336], bl[337], bl[338], bl[339], bl[340], bl[341], bl[342], bl[343], bl[344], bl[345], bl[346], bl[347], bl[348], bl[349], bl[350], bl[351], bl[352], bl[353], bl[354], bl[355], bl[356], bl[357], bl[358], bl[359], bl[360], bl[361], bl[362], bl[363], bl[364], bl[365], bl[366], bl[367], bl[368], bl[369], bl[370], bl[371], bl[372], bl[373], bl[374], bl[375], bl[17888], bl[17889], bl[17890], bl[17891], bl[17892], bl[17893], bl[17894], bl[17895], bl[17896], bl[17897], bl[17898], bl[17899], bl[17900], bl[17901], bl[17902], bl[17903], bl[17904], bl[17905], bl[17906], bl[17907], bl[17908], bl[17909], bl[17910], bl[17911], bl[17912], bl[17913], bl[17914], bl[17915], bl[17916], bl[17917], bl[17918], bl[17919], bl[17920], bl[17921], bl[17922], bl[17923], bl[17924], bl[17925], bl[17926], bl[17927], bl[17928], bl[17929], bl[17930], bl[17931], bl[17932], bl[17933], bl[17934], bl[17935], bl[17936], bl[17937], bl[17938], bl[17939], bl[17940], bl[17941], bl[17942], bl[17943], bl[17944], bl[17945], bl[17946], bl[17947], bl[17948], bl[17949], bl[17950], bl[17951], bl[17952], bl[17953], bl[17954], bl[17955], bl[17956], bl[17957], bl[17958], bl[17959], bl[17960], bl[17961], bl[17962], bl[17963], bl[17964], bl[17965], bl[17966], bl[17967], bl[224], bl[225], bl[226], bl[227], bl[228], bl[229], bl[230], bl[231], bl[232], bl[233], bl[234], bl[235], bl[236], bl[237], bl[238], bl[239], bl[240], bl[241], bl[242], bl[243], bl[244], bl[245], bl[246], bl[247], bl[248], bl[249], bl[250], bl[251], bl[252], bl[253], bl[254], bl[255], bl[256], bl[257], bl[258], bl[259], bl[260], bl[261], bl[262], bl[263], bl[264], bl[265], bl[266], bl[267], bl[268], bl[269], bl[270], bl[271], bl[272], bl[273], bl[274], bl[275], bl[276], bl[277], bl[278], bl[279], bl[280], bl[281], bl[282], bl[283], bl[284], bl[285], bl[286], bl[287], bl[288], bl[289], bl[290], bl[291], bl[292], bl[293], bl[294], bl[295], bl[296], bl[297], bl[298], bl[299], bl[300], bl[301], bl[302], bl[303]}),
        .wl({wl[17968], wl[17969], wl[17970], wl[17971], wl[17972], wl[17973], wl[17974], wl[17975], wl[17976], wl[17977], wl[17978], wl[17979], wl[17980], wl[17981], wl[17982], wl[17983], wl[17984], wl[17985], wl[17986], wl[17987], wl[17988], wl[17989], wl[17990], wl[17991], wl[17992], wl[17993], wl[17994], wl[17995], wl[17996], wl[17997], wl[17998], wl[17999], wl[18000], wl[18001], wl[18002], wl[18003], wl[18004], wl[18005], wl[18006], wl[18007], wl[18008], wl[18009], wl[18010], wl[18011], wl[18012], wl[18013], wl[18014], wl[18015], wl[18016], wl[18017], wl[18018], wl[18019], wl[18020], wl[18021], wl[18022], wl[18023], wl[18024], wl[18025], wl[18026], wl[18027], wl[18028], wl[18029], wl[18030], wl[18031], wl[18032], wl[18033], wl[18034], wl[18035], wl[18036], wl[18037], wl[18038], wl[18039], wl[18040], wl[18041], wl[18042], wl[18043], wl[18044], wl[18045], wl[18046], wl[18047], wl[18048], wl[18049], wl[18050], wl[18051], wl[18052], wl[18053], wl[18054], wl[18055], wl[18056], wl[18057], wl[18058], wl[18059], wl[18060], wl[18061], wl[18062], wl[18063], wl[18064], wl[18065], wl[18066], wl[18067], wl[18068], wl[18069], wl[18070], wl[18071], wl[18072], wl[18073], wl[18074], wl[18075], wl[18076], wl[18077], wl[18078], wl[18079], wl[18080], wl[18081], wl[18082], wl[18083], wl[18084], wl[18085], wl[18086], wl[18087], wl[18088], wl[18089], wl[18090], wl[18091], wl[18092], wl[18093], wl[18094], wl[18095], wl[18096], wl[18097], wl[18098], wl[18099], wl[18100], wl[18101], wl[18102], wl[18103], wl[18104], wl[18105], wl[18106], wl[18107], wl[18108], wl[18109], wl[18110], wl[18111], wl[18112], wl[18113], wl[18114], wl[18115], wl[18116], wl[18117], wl[18118], wl[18119], wl[18120], wl[18121], wl[18122], wl[18123], wl[18124], wl[18125], wl[18126], wl[18127], wl[18128], wl[18129], wl[18130], wl[18131], wl[18132], wl[18133], wl[18134], wl[18135], wl[18136], wl[18137], wl[18138], wl[18139], wl[18140], wl[18141], wl[18142], wl[18143], wl[18144], wl[18145], wl[18146], wl[18147], wl[18148], wl[18149], wl[18150], wl[18151], wl[18152], wl[18153], wl[18154], wl[18155], wl[18156], wl[18157], wl[18158], wl[18159], wl[18160], wl[18161], wl[18162], wl[18163], wl[18164], wl[18165], wl[18166], wl[18167], wl[18168], wl[18169], wl[18170], wl[18171], wl[18172], wl[18173], wl[18174], wl[18175], wl[18176], wl[18177], wl[18178], wl[18179], wl[18180], wl[18181], wl[18182], wl[18183], wl[18184], wl[18185], wl[18186], wl[18187], wl[18188], wl[18189], wl[18190], wl[18191], wl[18192], wl[18193], wl[18194], wl[18195], wl[18196], wl[18197], wl[18198], wl[18199], wl[18200], wl[18201], wl[18202], wl[18203], wl[18204], wl[18205], wl[18206], wl[18207], wl[18208], wl[18209], wl[18210], wl[18211], wl[18212], wl[18213], wl[18214], wl[18215], wl[18216], wl[18217], wl[18218], wl[18219], wl[18220], wl[18221], wl[18222], wl[18223], wl[18224], wl[18225], wl[18226], wl[18227], wl[18228], wl[18229], wl[18230], wl[18231], wl[18232], wl[18233], wl[18234], wl[18235], wl[18236], wl[18237], wl[18238], wl[18239], wl[18240], wl[18241], wl[18242], wl[18243], wl[18244], wl[18245], wl[18246], wl[18247], wl[18248], wl[18249], wl[18250], wl[18251], wl[18252], wl[18253], wl[18254], wl[18255], wl[18256], wl[18257], wl[18258], wl[18259], wl[18260], wl[18261], wl[18262], wl[18263], wl[18264], wl[18265], wl[18266], wl[18267], wl[18268], wl[18269], wl[18270], wl[18271], wl[18272], wl[18273], wl[18274], wl[18275], wl[18276], wl[18277], wl[18278], wl[18279], wl[18280], wl[18281], wl[18282], wl[18283], wl[18284], wl[18285], wl[18286], wl[18287], wl[18288], wl[18289], wl[18290], wl[18291], wl[18292], wl[18293], wl[18294], wl[18295], wl[18296], wl[18297], wl[18298], wl[18299], wl[18300], wl[18301], wl[18302], wl[18303], wl[18304], wl[18305], wl[18306], wl[18307], wl[18308], wl[18309], wl[18310], wl[18311], wl[18312], wl[18313], wl[18314], wl[18315], wl[18316], wl[18317], wl[18318], wl[18319], wl[18320], wl[18321], wl[18322], wl[18323], wl[18324], wl[18325], wl[18326], wl[18327], wl[18328], wl[18329], wl[18330], wl[18331], wl[18332], wl[18333], wl[18334], wl[18335], wl[18336], wl[18337], wl[18338], wl[18339], wl[18340], wl[18341], wl[18342], wl[18343], wl[18344], wl[18345], wl[18346], wl[18347], wl[18348], wl[18349], wl[18350], wl[18351], wl[18352], wl[18353], wl[18354], wl[18355], wl[18356], wl[18357], wl[18358], wl[18359], wl[18360], wl[18361], wl[18362], wl[18363], wl[18364], wl[18365], wl[18366], wl[18367], wl[18368], wl[18369], wl[18370], wl[18371], wl[18372], wl[18373], wl[18374], wl[18375], wl[18376], wl[18377], wl[18378], wl[18379], wl[18380], wl[18381], wl[18382], wl[18383], wl[18384], wl[18385], wl[18386], wl[18387], wl[18388], wl[18389], wl[18390], wl[18391], wl[18392], wl[18393], wl[18394], wl[18395], wl[18396], wl[18397], wl[18398], wl[18399], wl[18400], wl[18401], wl[18402], wl[18403], wl[18404], wl[18405], wl[18406], wl[18407], wl[18408], wl[18409], wl[18410], wl[18411], wl[18412], wl[18413], wl[18414], wl[18415], wl[18416], wl[18417], wl[18418], wl[18419], wl[18420], wl[18421], wl[18422], wl[18423], wl[18424], wl[18425], wl[18426], wl[18427], wl[18428], wl[18429], wl[18430], wl[18431], wl[18432], wl[18433], wl[18434], wl[18435], wl[18436], wl[18437], wl[18438], wl[18439], wl[18440], wl[18441], wl[18442], wl[18443], wl[18444], wl[18445], wl[18446], wl[18447], wl[18448], wl[18449], wl[18450], wl[18451], wl[18452], wl[18453], wl[18454], wl[18455], wl[18456], wl[18457], wl[18458], wl[18459], wl[18460], wl[18461], wl[18462], wl[18463], wl[18464], wl[18465], wl[18466], wl[18467], wl[18468], wl[18469], wl[18470], wl[18471], wl[18472], wl[18473], wl[18474], wl[18475], wl[18476], wl[18477], wl[18478], wl[18479], wl[18480], wl[18481], wl[18482], wl[18483], wl[18484], wl[18485], wl[18486], wl[18487], wl[18488], wl[18489], wl[18490], wl[18491], wl[18492], wl[18493], wl[18494], wl[18495], wl[18496], wl[18497], wl[18498], wl[18499], wl[18500], wl[18501], wl[18502], wl[18503], wl[18504], wl[18505], wl[18506], wl[18507], wl[18508], wl[18509], wl[18510], wl[18511], wl[18512], wl[18513], wl[18514], wl[18515], wl[18516], wl[18517], wl[18518], wl[18519], wl[18520], wl[18521], wl[18522], wl[18523], wl[18524], wl[18525], wl[18526], wl[18527], wl[18528], wl[18529], wl[18530], wl[18531], wl[18532], wl[18533], wl[18534], wl[18535], wl[18536], wl[18537], wl[18538], wl[18539], wl[18540], wl[18541], wl[18542], wl[18543], wl[18544], wl[18545], wl[18546], wl[18547], wl[18548], wl[18549], wl[18550], wl[18551], wl[18552], wl[18553], wl[18554], wl[18555], wl[18556], wl[18557], wl[18558], wl[18559], wl[18560], wl[18561], wl[18562], wl[18563], wl[18564], wl[18565], wl[18566], wl[18567], wl[18568], wl[18569], wl[18570], wl[18571], wl[18572], wl[18573], wl[18574], wl[18575], wl[18576], wl[18577], wl[18578], wl[18579], wl[18580], wl[18581], wl[18582], wl[18583], wl[18584], wl[18585], wl[18586], wl[18587], wl[18588], wl[18589], wl[18590], wl[18591], wl[18592], wl[18593], wl[18594], wl[18595], wl[18596], wl[18597], wl[18598], wl[18599], wl[18600], wl[18601], wl[18602], wl[18603], wl[18604], wl[18605], wl[18606], wl[18607], wl[18608], wl[18609], wl[18610], wl[18611], wl[18612], wl[18613], wl[18614], wl[18615], wl[18616], wl[18617], wl[18618], wl[18619], wl[18620], wl[18621], wl[18622], wl[18623], wl[18624], wl[18625], wl[18626], wl[18627], wl[18628], wl[18629], wl[18630], wl[18631], wl[18632], wl[18633], wl[18634], wl[18635], wl[18636], wl[18637], wl[18638], wl[18639], wl[18640], wl[18641], wl[18642], wl[18643], wl[18644], wl[18645], wl[18646], wl[18647], wl[18648], wl[18649], wl[18650], wl[18651], wl[18652], wl[18653], wl[18654], wl[18655], wl[18656], wl[18657], wl[18658], wl[18659], wl[18660], wl[18661], wl[18662], wl[18663], wl[18664], wl[18665], wl[18666], wl[18667], wl[18668], wl[18669], wl[18670], wl[18671], wl[18672], wl[18673], wl[18674], wl[18675], wl[18676], wl[18677], wl[18678], wl[18679], wl[18680], wl[18681], wl[18682], wl[18683], wl[18684], wl[18685], wl[18686], wl[18687], wl[18688], wl[18689], wl[18690], wl[18691], wl[18692], wl[18693], wl[18694], wl[18695], wl[18696], wl[18697], wl[18698], wl[18699], wl[18700], wl[18701], wl[18702], wl[18703], wl[18704], wl[18705], wl[18706], wl[18707], wl[18708], wl[18709], wl[18710], wl[18711], wl[18712], wl[18713], wl[18714], wl[18715], wl[18716], wl[18717], wl[18718], wl[18719], wl[18720], wl[18721], wl[18722], wl[18723], wl[18724], wl[18725], wl[18726], wl[18727], wl[18728], wl[18729], wl[18730], wl[18731], wl[18732], wl[18733], wl[18734], wl[18735], wl[18736], wl[18737], wl[18738], wl[18739], wl[18740], wl[18741], wl[18742], wl[18743], wl[18744], wl[18745], wl[18746], wl[18747], wl[18748], wl[18749], wl[18750], wl[18751], wl[18752], wl[18753], wl[18754], wl[18755], wl[18756], wl[18757], wl[18758], wl[18759], wl[18760], wl[18761], wl[18762], wl[18763], wl[18764], wl[18765], wl[18766], wl[18767], wl[18768], wl[18769], wl[18770], wl[18771], wl[18772], wl[18773], wl[18774], wl[18775], wl[18776], wl[18777], wl[18778], wl[18779], wl[18780], wl[18781], wl[18782], wl[18783], wl[18784], wl[18785], wl[18786], wl[18787], wl[18788], wl[18789], wl[18790], wl[18791], wl[18792], wl[18793], wl[18794], wl[18795], wl[18796], wl[18797], wl[18798], wl[18799], wl[18800], wl[18801], wl[18802], wl[18803], wl[18804], wl[18805], wl[18806], wl[18807], wl[18808], wl[18809], wl[18810], wl[18811], wl[18812], wl[18813], wl[18814], wl[18815], wl[18816], wl[18817], wl[18818], wl[18819], wl[18820], wl[18821], wl[18822], wl[18823], wl[18824], wl[18825], wl[18826], wl[18827], wl[18828], wl[18829], wl[18830], wl[18831], wl[18832], wl[18833], wl[18834], wl[18835], wl[18836], wl[18837], wl[18838], wl[18839], wl[18840], wl[18841], wl[18842], wl[18843], wl[18844], wl[18845], wl[18846], wl[18847], wl[18848], wl[18849], wl[18850], wl[18851], wl[18852], wl[18853], wl[18854], wl[18855], wl[18856], wl[18857], wl[18858], wl[18859], wl[18860], wl[18861], wl[18862], wl[18863], wl[18864], wl[18865], wl[18866], wl[18867], wl[18868], wl[18869], wl[18870], wl[18871], wl[18872], wl[18873], wl[18874], wl[18875], wl[18876], wl[18877], wl[18878], wl[18879], wl[18880], wl[18881], wl[18882], wl[18883], wl[18884], wl[18885], wl[18886], wl[18887], wl[18888], wl[18889], wl[18890], wl[18891], wl[18892], wl[18893], wl[18894], wl[18895], wl[18896], wl[18897], wl[18898], wl[18899], wl[18900], wl[18901], wl[18902], wl[18903], wl[18904], wl[18905], wl[18906], wl[18907], wl[18908], wl[18909], wl[18910], wl[18911], wl[18912], wl[18913], wl[18914], wl[18915], wl[18916], wl[18917], wl[18918], wl[18919], wl[18920], wl[18921], wl[18922], wl[18923], wl[18924], wl[18925], wl[18926], wl[18927], wl[18928], wl[18929], wl[18930], wl[18931], wl[18932], wl[18933], wl[18934], wl[18935], wl[18936], wl[18937], wl[18938], wl[18939], wl[18940], wl[18941], wl[18942], wl[18943], wl[18944], wl[18945], wl[18946], wl[18947], wl[18948], wl[18949], wl[18950], wl[18951], wl[18952], wl[18953], wl[18954], wl[18955], wl[18956], wl[18957], wl[18958], wl[18959], wl[18960], wl[18961], wl[18962], wl[18963], wl[18964], wl[18965], wl[18966], wl[18967], wl[18968], wl[18969], wl[18970], wl[18971], wl[18972], wl[18973], wl[18974], wl[18975], wl[18976], wl[18977], wl[18978], wl[18979], wl[18980], wl[18981], wl[18982], wl[18983], wl[18984], wl[18985], wl[18986], wl[18987], wl[376], wl[377], wl[378], wl[379], wl[380], wl[381], wl[382], wl[383], wl[304], wl[305], wl[306], wl[307], wl[308], wl[309], wl[310], wl[311], wl[312], wl[313], wl[314], wl[315], wl[316], wl[317], wl[318], wl[319], wl[320], wl[321], wl[322], wl[323], wl[324], wl[325], wl[326], wl[327], wl[328], wl[329], wl[330], wl[331], wl[332], wl[333], wl[334], wl[335], wl[336], wl[337], wl[338], wl[339], wl[340], wl[341], wl[342], wl[343], wl[344], wl[345], wl[346], wl[347], wl[348], wl[349], wl[350], wl[351], wl[352], wl[353], wl[354], wl[355], wl[356], wl[357], wl[358], wl[359], wl[360], wl[361], wl[362], wl[363], wl[364], wl[365], wl[366], wl[367], wl[368], wl[369], wl[370], wl[371], wl[372], wl[373], wl[374], wl[375], wl[17888], wl[17889], wl[17890], wl[17891], wl[17892], wl[17893], wl[17894], wl[17895], wl[17896], wl[17897], wl[17898], wl[17899], wl[17900], wl[17901], wl[17902], wl[17903], wl[17904], wl[17905], wl[17906], wl[17907], wl[17908], wl[17909], wl[17910], wl[17911], wl[17912], wl[17913], wl[17914], wl[17915], wl[17916], wl[17917], wl[17918], wl[17919], wl[17920], wl[17921], wl[17922], wl[17923], wl[17924], wl[17925], wl[17926], wl[17927], wl[17928], wl[17929], wl[17930], wl[17931], wl[17932], wl[17933], wl[17934], wl[17935], wl[17936], wl[17937], wl[17938], wl[17939], wl[17940], wl[17941], wl[17942], wl[17943], wl[17944], wl[17945], wl[17946], wl[17947], wl[17948], wl[17949], wl[17950], wl[17951], wl[17952], wl[17953], wl[17954], wl[17955], wl[17956], wl[17957], wl[17958], wl[17959], wl[17960], wl[17961], wl[17962], wl[17963], wl[17964], wl[17965], wl[17966], wl[17967], wl[224], wl[225], wl[226], wl[227], wl[228], wl[229], wl[230], wl[231], wl[232], wl[233], wl[234], wl[235], wl[236], wl[237], wl[238], wl[239], wl[240], wl[241], wl[242], wl[243], wl[244], wl[245], wl[246], wl[247], wl[248], wl[249], wl[250], wl[251], wl[252], wl[253], wl[254], wl[255], wl[256], wl[257], wl[258], wl[259], wl[260], wl[261], wl[262], wl[263], wl[264], wl[265], wl[266], wl[267], wl[268], wl[269], wl[270], wl[271], wl[272], wl[273], wl[274], wl[275], wl[276], wl[277], wl[278], wl[279], wl[280], wl[281], wl[282], wl[283], wl[284], wl[285], wl[286], wl[287], wl[288], wl[289], wl[290], wl[291], wl[292], wl[293], wl[294], wl[295], wl[296], wl[297], wl[298], wl[299], wl[300], wl[301], wl[302], wl[303]})
    );
    top_left_tile tile_1__5_
    (
        .chanx_right_in(cbx_1__4__0_chanx_left_out),
        .chanx_right_out(sb_0__4__0_chanx_right_out),
        .grid_right_t_inpad(grid_io_top_1__5__io_bottom_in),
        .grid_right_b_in(sb_0__4__grid_right_b_in),
        .grid_bottom_r_in(sb_0__3__grid_top_r_in),
        .grid_bottom_l_inpad(grid_io_left_0__4__io_right_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[120:127]),
        .chany_bottom_in_0(sb_0__1__2_chany_top_out),
        .chany_bottom_out_0(cby_0__1__3_chany_bottom_out),
        .grid_right_out(grid_clb_1__4__grid_left_in),
        .bl({bl[704], bl[705], bl[706], bl[707], bl[708], bl[709], bl[710], bl[711], bl[712], bl[713], bl[714], bl[715], bl[716], bl[717], bl[718], bl[719], bl[720], bl[721], bl[722], bl[723], bl[724], bl[725], bl[726], bl[727], bl[728], bl[729], bl[730], bl[731], bl[732], bl[733], bl[734], bl[735], bl[736], bl[737], bl[738], bl[739], bl[740], bl[741], bl[742], bl[743], bl[744], bl[745], bl[746], bl[747], bl[748], bl[749], bl[750], bl[751], bl[752], bl[753], bl[754], bl[755], bl[756], bl[757], bl[758], bl[759], bl[760], bl[761], bl[762], bl[763], bl[764], bl[765], bl[766], bl[767], bl[768], bl[769], bl[770], bl[771], bl[772], bl[773], bl[774], bl[775], bl[776], bl[777], bl[778], bl[779], bl[780], bl[781], bl[782], bl[783], bl[934], bl[935], bl[936], bl[937], bl[938], bl[939], bl[940], bl[941], bl[862], bl[863], bl[864], bl[865], bl[866], bl[867], bl[868], bl[869], bl[870], bl[871], bl[872], bl[873], bl[874], bl[875], bl[876], bl[877], bl[878], bl[879], bl[880], bl[881], bl[882], bl[883], bl[884], bl[885], bl[886], bl[887], bl[888], bl[889], bl[890], bl[891], bl[892], bl[893], bl[894], bl[895], bl[896], bl[897], bl[898], bl[899], bl[900], bl[901], bl[902], bl[903], bl[904], bl[905], bl[906], bl[907], bl[908], bl[909], bl[910], bl[911], bl[912], bl[913], bl[914], bl[915], bl[916], bl[917], bl[918], bl[919], bl[920], bl[921], bl[922], bl[923], bl[924], bl[925], bl[926], bl[927], bl[928], bl[929], bl[930], bl[931], bl[932], bl[933]}),
        .wl({wl[704], wl[705], wl[706], wl[707], wl[708], wl[709], wl[710], wl[711], wl[712], wl[713], wl[714], wl[715], wl[716], wl[717], wl[718], wl[719], wl[720], wl[721], wl[722], wl[723], wl[724], wl[725], wl[726], wl[727], wl[728], wl[729], wl[730], wl[731], wl[732], wl[733], wl[734], wl[735], wl[736], wl[737], wl[738], wl[739], wl[740], wl[741], wl[742], wl[743], wl[744], wl[745], wl[746], wl[747], wl[748], wl[749], wl[750], wl[751], wl[752], wl[753], wl[754], wl[755], wl[756], wl[757], wl[758], wl[759], wl[760], wl[761], wl[762], wl[763], wl[764], wl[765], wl[766], wl[767], wl[768], wl[769], wl[770], wl[771], wl[772], wl[773], wl[774], wl[775], wl[776], wl[777], wl[778], wl[779], wl[780], wl[781], wl[782], wl[783], wl[934], wl[935], wl[936], wl[937], wl[938], wl[939], wl[940], wl[941], wl[862], wl[863], wl[864], wl[865], wl[866], wl[867], wl[868], wl[869], wl[870], wl[871], wl[872], wl[873], wl[874], wl[875], wl[876], wl[877], wl[878], wl[879], wl[880], wl[881], wl[882], wl[883], wl[884], wl[885], wl[886], wl[887], wl[888], wl[889], wl[890], wl[891], wl[892], wl[893], wl[894], wl[895], wl[896], wl[897], wl[898], wl[899], wl[900], wl[901], wl[902], wl[903], wl[904], wl[905], wl[906], wl[907], wl[908], wl[909], wl[910], wl[911], wl[912], wl[913], wl[914], wl[915], wl[916], wl[917], wl[918], wl[919], wl[920], wl[921], wl[922], wl[923], wl[924], wl[925], wl[926], wl[927], wl[928], wl[929], wl[930], wl[931], wl[932], wl[933]})
    );
    top_right_tile tile_5__5_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_3__4__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_3__4__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_3__4__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_4__3__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_4__3__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_4__3__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_3__3__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_3__3__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_3__3__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_3__3__grid_top_r_in[1]),
        .grid_left_in(grid_clb_4__4__grid_left_in),
        .grid_bottom_in(grid_clb_4__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[24:31]),
        .io_bottom_in(grid_io_top_4__5__io_bottom_in),
        .chanx_left_in(sb_1__4__2_chanx_right_out),
        .chanx_left_out(cbx_1__4__3_chanx_left_out),
        .gfpga_pad_GPIO_PAD_0(gfpga_pad_GPIO_PAD[32:39]),
        .io_left_in(grid_io_right_5__4__io_left_in),
        .chany_bottom_in(sb_4__1__2_chany_top_out),
        .chany_bottom_out(cby_4__1__3_chany_bottom_out),
        .grid_bottom_l_in(sb_4__3__grid_top_l_in),
        .grid_left_b_in(sb_3__4__grid_right_b_in),
        .bl({bl[16708], bl[16709], bl[16710], bl[16711], bl[16712], bl[16713], bl[16714], bl[16715], bl[16716], bl[16717], bl[16718], bl[16719], bl[16720], bl[16721], bl[16722], bl[16723], bl[16724], bl[16725], bl[16726], bl[16727], bl[16728], bl[16729], bl[16730], bl[16731], bl[16732], bl[16733], bl[16734], bl[16735], bl[16736], bl[16737], bl[16738], bl[16739], bl[16740], bl[16741], bl[16742], bl[16743], bl[16744], bl[16745], bl[16746], bl[16747], bl[16748], bl[16749], bl[16750], bl[16751], bl[16752], bl[16753], bl[16754], bl[16755], bl[16756], bl[16757], bl[16758], bl[16759], bl[16760], bl[16761], bl[16762], bl[16763], bl[16764], bl[16765], bl[16766], bl[16767], bl[16768], bl[16769], bl[16770], bl[16771], bl[16772], bl[16773], bl[16774], bl[16775], bl[16776], bl[16777], bl[16778], bl[16779], bl[16780], bl[16781], bl[16782], bl[16783], bl[16784], bl[16785], bl[16786], bl[16787], bl[16788], bl[16789], bl[16790], bl[16791], bl[16792], bl[16793], bl[16794], bl[16795], bl[16796], bl[16797], bl[16798], bl[16799], bl[16800], bl[16801], bl[16802], bl[16803], bl[16804], bl[16805], bl[16806], bl[16807], bl[16808], bl[16809], bl[16810], bl[16811], bl[16812], bl[16813], bl[16814], bl[16815], bl[16816], bl[16817], bl[16818], bl[16819], bl[16820], bl[16821], bl[16822], bl[16823], bl[16824], bl[16825], bl[16826], bl[16827], bl[16828], bl[16829], bl[16830], bl[16831], bl[16832], bl[16833], bl[16834], bl[16835], bl[16836], bl[16837], bl[16838], bl[16839], bl[16840], bl[16841], bl[16842], bl[16843], bl[16844], bl[16845], bl[16846], bl[16847], bl[16848], bl[16849], bl[16850], bl[16851], bl[16852], bl[16853], bl[16854], bl[16855], bl[16856], bl[16857], bl[16858], bl[16859], bl[16860], bl[16861], bl[16862], bl[16863], bl[16864], bl[16865], bl[16866], bl[16867], bl[16868], bl[16869], bl[16870], bl[16871], bl[16872], bl[16873], bl[16874], bl[16875], bl[16876], bl[16877], bl[16878], bl[16879], bl[16880], bl[16881], bl[16882], bl[16883], bl[16884], bl[16885], bl[16886], bl[16887], bl[16888], bl[16889], bl[16890], bl[16891], bl[16892], bl[16893], bl[16894], bl[16895], bl[16896], bl[16897], bl[16898], bl[16899], bl[16900], bl[16901], bl[16902], bl[16903], bl[16904], bl[16905], bl[16906], bl[16907], bl[16908], bl[16909], bl[16910], bl[16911], bl[16912], bl[16913], bl[16914], bl[16915], bl[16916], bl[16917], bl[16918], bl[16919], bl[16920], bl[16921], bl[16922], bl[16923], bl[16924], bl[16925], bl[16926], bl[16927], bl[16928], bl[16929], bl[16930], bl[16931], bl[16932], bl[16933], bl[16934], bl[16935], bl[16936], bl[16937], bl[16938], bl[16939], bl[16940], bl[16941], bl[16942], bl[16943], bl[16944], bl[16945], bl[16946], bl[16947], bl[16948], bl[16949], bl[16950], bl[16951], bl[16952], bl[16953], bl[16954], bl[16955], bl[16956], bl[16957], bl[16958], bl[16959], bl[16960], bl[16961], bl[16962], bl[16963], bl[16964], bl[16965], bl[16966], bl[16967], bl[16968], bl[16969], bl[16970], bl[16971], bl[16972], bl[16973], bl[16974], bl[16975], bl[16976], bl[16977], bl[16978], bl[16979], bl[16980], bl[16981], bl[16982], bl[16983], bl[16984], bl[16985], bl[16986], bl[16987], bl[16988], bl[16989], bl[16990], bl[16991], bl[16992], bl[16993], bl[16994], bl[16995], bl[16996], bl[16997], bl[16998], bl[16999], bl[17000], bl[17001], bl[17002], bl[17003], bl[17004], bl[17005], bl[17006], bl[17007], bl[17008], bl[17009], bl[17010], bl[17011], bl[17012], bl[17013], bl[17014], bl[17015], bl[17016], bl[17017], bl[17018], bl[17019], bl[17020], bl[17021], bl[17022], bl[17023], bl[17024], bl[17025], bl[17026], bl[17027], bl[17028], bl[17029], bl[17030], bl[17031], bl[17032], bl[17033], bl[17034], bl[17035], bl[17036], bl[17037], bl[17038], bl[17039], bl[17040], bl[17041], bl[17042], bl[17043], bl[17044], bl[17045], bl[17046], bl[17047], bl[17048], bl[17049], bl[17050], bl[17051], bl[17052], bl[17053], bl[17054], bl[17055], bl[17056], bl[17057], bl[17058], bl[17059], bl[17060], bl[17061], bl[17062], bl[17063], bl[17064], bl[17065], bl[17066], bl[17067], bl[17068], bl[17069], bl[17070], bl[17071], bl[17072], bl[17073], bl[17074], bl[17075], bl[17076], bl[17077], bl[17078], bl[17079], bl[17080], bl[17081], bl[17082], bl[17083], bl[17084], bl[17085], bl[17086], bl[17087], bl[17088], bl[17089], bl[17090], bl[17091], bl[17092], bl[17093], bl[17094], bl[17095], bl[17096], bl[17097], bl[17098], bl[17099], bl[17100], bl[17101], bl[17102], bl[17103], bl[17104], bl[17105], bl[17106], bl[17107], bl[17108], bl[17109], bl[17110], bl[17111], bl[17112], bl[17113], bl[17114], bl[17115], bl[17116], bl[17117], bl[17118], bl[17119], bl[17120], bl[17121], bl[17122], bl[17123], bl[17124], bl[17125], bl[17126], bl[17127], bl[17128], bl[17129], bl[17130], bl[17131], bl[17132], bl[17133], bl[17134], bl[17135], bl[17136], bl[17137], bl[17138], bl[17139], bl[17140], bl[17141], bl[17142], bl[17143], bl[17144], bl[17145], bl[17146], bl[17147], bl[17148], bl[17149], bl[17150], bl[17151], bl[17152], bl[17153], bl[17154], bl[17155], bl[17156], bl[17157], bl[17158], bl[17159], bl[17160], bl[17161], bl[17162], bl[17163], bl[17164], bl[17165], bl[17166], bl[17167], bl[17168], bl[17169], bl[17170], bl[17171], bl[17172], bl[17173], bl[17174], bl[17175], bl[17176], bl[17177], bl[17178], bl[17179], bl[17180], bl[17181], bl[17182], bl[17183], bl[17184], bl[17185], bl[17186], bl[17187], bl[17188], bl[17189], bl[17190], bl[17191], bl[17192], bl[17193], bl[17194], bl[17195], bl[17196], bl[17197], bl[17198], bl[17199], bl[17200], bl[17201], bl[17202], bl[17203], bl[17204], bl[17205], bl[17206], bl[17207], bl[17208], bl[17209], bl[17210], bl[17211], bl[17212], bl[17213], bl[17214], bl[17215], bl[17216], bl[17217], bl[17218], bl[17219], bl[17220], bl[17221], bl[17222], bl[17223], bl[17224], bl[17225], bl[17226], bl[17227], bl[17228], bl[17229], bl[17230], bl[17231], bl[17232], bl[17233], bl[17234], bl[17235], bl[17236], bl[17237], bl[17238], bl[17239], bl[17240], bl[17241], bl[17242], bl[17243], bl[17244], bl[17245], bl[17246], bl[17247], bl[17248], bl[17249], bl[17250], bl[17251], bl[17252], bl[17253], bl[17254], bl[17255], bl[17256], bl[17257], bl[17258], bl[17259], bl[17260], bl[17261], bl[17262], bl[17263], bl[17264], bl[17265], bl[17266], bl[17267], bl[17268], bl[17269], bl[17270], bl[17271], bl[17272], bl[17273], bl[17274], bl[17275], bl[17276], bl[17277], bl[17278], bl[17279], bl[17280], bl[17281], bl[17282], bl[17283], bl[17284], bl[17285], bl[17286], bl[17287], bl[17288], bl[17289], bl[17290], bl[17291], bl[17292], bl[17293], bl[17294], bl[17295], bl[17296], bl[17297], bl[17298], bl[17299], bl[17300], bl[17301], bl[17302], bl[17303], bl[17304], bl[17305], bl[17306], bl[17307], bl[17308], bl[17309], bl[17310], bl[17311], bl[17312], bl[17313], bl[17314], bl[17315], bl[17316], bl[17317], bl[17318], bl[17319], bl[17320], bl[17321], bl[17322], bl[17323], bl[17324], bl[17325], bl[17326], bl[17327], bl[17328], bl[17329], bl[17330], bl[17331], bl[17332], bl[17333], bl[17334], bl[17335], bl[17336], bl[17337], bl[17338], bl[17339], bl[17340], bl[17341], bl[17342], bl[17343], bl[17344], bl[17345], bl[17346], bl[17347], bl[17348], bl[17349], bl[17350], bl[17351], bl[17352], bl[17353], bl[17354], bl[17355], bl[17356], bl[17357], bl[17358], bl[17359], bl[17360], bl[17361], bl[17362], bl[17363], bl[17364], bl[17365], bl[17366], bl[17367], bl[17368], bl[17369], bl[17370], bl[17371], bl[17372], bl[17373], bl[17374], bl[17375], bl[17376], bl[17377], bl[17378], bl[17379], bl[17380], bl[17381], bl[17382], bl[17383], bl[17384], bl[17385], bl[17386], bl[17387], bl[17388], bl[17389], bl[17390], bl[17391], bl[17392], bl[17393], bl[17394], bl[17395], bl[17396], bl[17397], bl[17398], bl[17399], bl[17400], bl[17401], bl[17402], bl[17403], bl[17404], bl[17405], bl[17406], bl[17407], bl[17408], bl[17409], bl[17410], bl[17411], bl[17412], bl[17413], bl[17414], bl[17415], bl[17416], bl[17417], bl[17418], bl[17419], bl[17420], bl[17421], bl[17422], bl[17423], bl[17424], bl[17425], bl[17426], bl[17427], bl[17428], bl[17429], bl[17430], bl[17431], bl[17432], bl[17433], bl[17434], bl[17435], bl[17436], bl[17437], bl[17438], bl[17439], bl[17440], bl[17441], bl[17442], bl[17443], bl[17444], bl[17445], bl[17446], bl[17447], bl[17448], bl[17449], bl[17450], bl[17451], bl[17452], bl[17453], bl[17454], bl[17455], bl[17456], bl[17457], bl[17458], bl[17459], bl[17460], bl[17461], bl[17462], bl[17463], bl[17464], bl[17465], bl[17466], bl[17467], bl[17468], bl[17469], bl[17470], bl[17471], bl[17472], bl[17473], bl[17474], bl[17475], bl[17476], bl[17477], bl[17478], bl[17479], bl[17480], bl[17481], bl[17482], bl[17483], bl[17484], bl[17485], bl[17486], bl[17487], bl[17488], bl[17489], bl[17490], bl[17491], bl[17492], bl[17493], bl[17494], bl[17495], bl[17496], bl[17497], bl[17498], bl[17499], bl[17500], bl[17501], bl[17502], bl[17503], bl[17504], bl[17505], bl[17506], bl[17507], bl[17508], bl[17509], bl[17510], bl[17511], bl[17512], bl[17513], bl[17514], bl[17515], bl[17516], bl[17517], bl[17518], bl[17519], bl[17520], bl[17521], bl[17522], bl[17523], bl[17524], bl[17525], bl[17526], bl[17527], bl[17528], bl[17529], bl[17530], bl[17531], bl[17532], bl[17533], bl[17534], bl[17535], bl[17536], bl[17537], bl[17538], bl[17539], bl[17540], bl[17541], bl[17542], bl[17543], bl[17544], bl[17545], bl[17546], bl[17547], bl[17548], bl[17549], bl[17550], bl[17551], bl[17552], bl[17553], bl[17554], bl[17555], bl[17556], bl[17557], bl[17558], bl[17559], bl[17560], bl[17561], bl[17562], bl[17563], bl[17564], bl[17565], bl[17566], bl[17567], bl[17568], bl[17569], bl[17570], bl[17571], bl[17572], bl[17573], bl[17574], bl[17575], bl[17576], bl[17577], bl[17578], bl[17579], bl[17580], bl[17581], bl[17582], bl[17583], bl[17584], bl[17585], bl[17586], bl[17587], bl[17588], bl[17589], bl[17590], bl[17591], bl[17592], bl[17593], bl[17594], bl[17595], bl[17596], bl[17597], bl[17598], bl[17599], bl[17600], bl[17601], bl[17602], bl[17603], bl[17604], bl[17605], bl[17606], bl[17607], bl[17608], bl[17609], bl[17610], bl[17611], bl[17612], bl[17613], bl[17614], bl[17615], bl[17616], bl[17617], bl[17618], bl[17619], bl[17620], bl[17621], bl[17622], bl[17623], bl[17624], bl[17625], bl[17626], bl[17627], bl[17628], bl[17629], bl[17630], bl[17631], bl[17632], bl[17633], bl[17634], bl[17635], bl[17636], bl[17637], bl[17638], bl[17639], bl[17640], bl[17641], bl[17642], bl[17643], bl[17644], bl[17645], bl[17646], bl[17647], bl[17648], bl[17649], bl[17650], bl[17651], bl[17652], bl[17653], bl[17654], bl[17655], bl[17656], bl[17657], bl[17658], bl[17659], bl[17660], bl[17661], bl[17662], bl[17663], bl[17664], bl[17665], bl[17666], bl[17667], bl[17668], bl[17669], bl[17670], bl[17671], bl[17672], bl[17673], bl[17674], bl[17675], bl[17676], bl[17677], bl[17678], bl[17679], bl[17680], bl[17681], bl[17682], bl[17683], bl[17684], bl[17685], bl[17686], bl[17687], bl[17688], bl[17689], bl[17690], bl[17691], bl[17692], bl[17693], bl[17694], bl[17695], bl[17696], bl[17697], bl[17698], bl[17699], bl[17700], bl[17701], bl[17702], bl[17703], bl[17704], bl[17705], bl[17706], bl[17707], bl[17708], bl[17709], bl[17710], bl[17711], bl[17712], bl[17713], bl[17714], bl[17715], bl[17716], bl[17717], bl[17718], bl[17719], bl[17720], bl[17721], bl[17722], bl[17723], bl[17724], bl[17725], bl[17726], bl[17727], bl[216], bl[217], bl[218], bl[219], bl[220], bl[221], bl[222], bl[223], bl[144], bl[145], bl[146], bl[147], bl[148], bl[149], bl[150], bl[151], bl[152], bl[153], bl[154], bl[155], bl[156], bl[157], bl[158], bl[159], bl[160], bl[161], bl[162], bl[163], bl[164], bl[165], bl[166], bl[167], bl[168], bl[169], bl[170], bl[171], bl[172], bl[173], bl[174], bl[175], bl[176], bl[177], bl[178], bl[179], bl[180], bl[181], bl[182], bl[183], bl[184], bl[185], bl[186], bl[187], bl[188], bl[189], bl[190], bl[191], bl[192], bl[193], bl[194], bl[195], bl[196], bl[197], bl[198], bl[199], bl[200], bl[201], bl[202], bl[203], bl[204], bl[205], bl[206], bl[207], bl[208], bl[209], bl[210], bl[211], bl[212], bl[213], bl[214], bl[215], bl[56], bl[57], bl[58], bl[59], bl[60], bl[61], bl[62], bl[63], bl[16636], bl[16637], bl[16638], bl[16639], bl[16640], bl[16641], bl[16642], bl[16643], bl[16644], bl[16645], bl[16646], bl[16647], bl[16648], bl[16649], bl[16650], bl[16651], bl[16652], bl[16653], bl[16654], bl[16655], bl[16656], bl[16657], bl[16658], bl[16659], bl[16660], bl[16661], bl[16662], bl[16663], bl[16664], bl[16665], bl[16666], bl[16667], bl[16668], bl[16669], bl[16670], bl[16671], bl[16672], bl[16673], bl[16674], bl[16675], bl[16676], bl[16677], bl[16678], bl[16679], bl[16680], bl[16681], bl[16682], bl[16683], bl[16684], bl[16685], bl[16686], bl[16687], bl[16688], bl[16689], bl[16690], bl[16691], bl[16692], bl[16693], bl[16694], bl[16695], bl[16696], bl[16697], bl[16698], bl[16699], bl[16700], bl[16701], bl[16702], bl[16703], bl[16704], bl[16705], bl[16706], bl[16707], bl[64], bl[65], bl[66], bl[67], bl[68], bl[69], bl[70], bl[71], bl[72], bl[73], bl[74], bl[75], bl[76], bl[77], bl[78], bl[79], bl[80], bl[81], bl[82], bl[83], bl[84], bl[85], bl[86], bl[87], bl[88], bl[89], bl[90], bl[91], bl[92], bl[93], bl[94], bl[95], bl[96], bl[97], bl[98], bl[99], bl[100], bl[101], bl[102], bl[103], bl[104], bl[105], bl[106], bl[107], bl[108], bl[109], bl[110], bl[111], bl[112], bl[113], bl[114], bl[115], bl[116], bl[117], bl[118], bl[119], bl[120], bl[121], bl[122], bl[123], bl[124], bl[125], bl[126], bl[127], bl[128], bl[129], bl[130], bl[131], bl[132], bl[133], bl[134], bl[135], bl[136], bl[137], bl[138], bl[139], bl[140], bl[141], bl[142], bl[143]}),
        .wl({wl[16708], wl[16709], wl[16710], wl[16711], wl[16712], wl[16713], wl[16714], wl[16715], wl[16716], wl[16717], wl[16718], wl[16719], wl[16720], wl[16721], wl[16722], wl[16723], wl[16724], wl[16725], wl[16726], wl[16727], wl[16728], wl[16729], wl[16730], wl[16731], wl[16732], wl[16733], wl[16734], wl[16735], wl[16736], wl[16737], wl[16738], wl[16739], wl[16740], wl[16741], wl[16742], wl[16743], wl[16744], wl[16745], wl[16746], wl[16747], wl[16748], wl[16749], wl[16750], wl[16751], wl[16752], wl[16753], wl[16754], wl[16755], wl[16756], wl[16757], wl[16758], wl[16759], wl[16760], wl[16761], wl[16762], wl[16763], wl[16764], wl[16765], wl[16766], wl[16767], wl[16768], wl[16769], wl[16770], wl[16771], wl[16772], wl[16773], wl[16774], wl[16775], wl[16776], wl[16777], wl[16778], wl[16779], wl[16780], wl[16781], wl[16782], wl[16783], wl[16784], wl[16785], wl[16786], wl[16787], wl[16788], wl[16789], wl[16790], wl[16791], wl[16792], wl[16793], wl[16794], wl[16795], wl[16796], wl[16797], wl[16798], wl[16799], wl[16800], wl[16801], wl[16802], wl[16803], wl[16804], wl[16805], wl[16806], wl[16807], wl[16808], wl[16809], wl[16810], wl[16811], wl[16812], wl[16813], wl[16814], wl[16815], wl[16816], wl[16817], wl[16818], wl[16819], wl[16820], wl[16821], wl[16822], wl[16823], wl[16824], wl[16825], wl[16826], wl[16827], wl[16828], wl[16829], wl[16830], wl[16831], wl[16832], wl[16833], wl[16834], wl[16835], wl[16836], wl[16837], wl[16838], wl[16839], wl[16840], wl[16841], wl[16842], wl[16843], wl[16844], wl[16845], wl[16846], wl[16847], wl[16848], wl[16849], wl[16850], wl[16851], wl[16852], wl[16853], wl[16854], wl[16855], wl[16856], wl[16857], wl[16858], wl[16859], wl[16860], wl[16861], wl[16862], wl[16863], wl[16864], wl[16865], wl[16866], wl[16867], wl[16868], wl[16869], wl[16870], wl[16871], wl[16872], wl[16873], wl[16874], wl[16875], wl[16876], wl[16877], wl[16878], wl[16879], wl[16880], wl[16881], wl[16882], wl[16883], wl[16884], wl[16885], wl[16886], wl[16887], wl[16888], wl[16889], wl[16890], wl[16891], wl[16892], wl[16893], wl[16894], wl[16895], wl[16896], wl[16897], wl[16898], wl[16899], wl[16900], wl[16901], wl[16902], wl[16903], wl[16904], wl[16905], wl[16906], wl[16907], wl[16908], wl[16909], wl[16910], wl[16911], wl[16912], wl[16913], wl[16914], wl[16915], wl[16916], wl[16917], wl[16918], wl[16919], wl[16920], wl[16921], wl[16922], wl[16923], wl[16924], wl[16925], wl[16926], wl[16927], wl[16928], wl[16929], wl[16930], wl[16931], wl[16932], wl[16933], wl[16934], wl[16935], wl[16936], wl[16937], wl[16938], wl[16939], wl[16940], wl[16941], wl[16942], wl[16943], wl[16944], wl[16945], wl[16946], wl[16947], wl[16948], wl[16949], wl[16950], wl[16951], wl[16952], wl[16953], wl[16954], wl[16955], wl[16956], wl[16957], wl[16958], wl[16959], wl[16960], wl[16961], wl[16962], wl[16963], wl[16964], wl[16965], wl[16966], wl[16967], wl[16968], wl[16969], wl[16970], wl[16971], wl[16972], wl[16973], wl[16974], wl[16975], wl[16976], wl[16977], wl[16978], wl[16979], wl[16980], wl[16981], wl[16982], wl[16983], wl[16984], wl[16985], wl[16986], wl[16987], wl[16988], wl[16989], wl[16990], wl[16991], wl[16992], wl[16993], wl[16994], wl[16995], wl[16996], wl[16997], wl[16998], wl[16999], wl[17000], wl[17001], wl[17002], wl[17003], wl[17004], wl[17005], wl[17006], wl[17007], wl[17008], wl[17009], wl[17010], wl[17011], wl[17012], wl[17013], wl[17014], wl[17015], wl[17016], wl[17017], wl[17018], wl[17019], wl[17020], wl[17021], wl[17022], wl[17023], wl[17024], wl[17025], wl[17026], wl[17027], wl[17028], wl[17029], wl[17030], wl[17031], wl[17032], wl[17033], wl[17034], wl[17035], wl[17036], wl[17037], wl[17038], wl[17039], wl[17040], wl[17041], wl[17042], wl[17043], wl[17044], wl[17045], wl[17046], wl[17047], wl[17048], wl[17049], wl[17050], wl[17051], wl[17052], wl[17053], wl[17054], wl[17055], wl[17056], wl[17057], wl[17058], wl[17059], wl[17060], wl[17061], wl[17062], wl[17063], wl[17064], wl[17065], wl[17066], wl[17067], wl[17068], wl[17069], wl[17070], wl[17071], wl[17072], wl[17073], wl[17074], wl[17075], wl[17076], wl[17077], wl[17078], wl[17079], wl[17080], wl[17081], wl[17082], wl[17083], wl[17084], wl[17085], wl[17086], wl[17087], wl[17088], wl[17089], wl[17090], wl[17091], wl[17092], wl[17093], wl[17094], wl[17095], wl[17096], wl[17097], wl[17098], wl[17099], wl[17100], wl[17101], wl[17102], wl[17103], wl[17104], wl[17105], wl[17106], wl[17107], wl[17108], wl[17109], wl[17110], wl[17111], wl[17112], wl[17113], wl[17114], wl[17115], wl[17116], wl[17117], wl[17118], wl[17119], wl[17120], wl[17121], wl[17122], wl[17123], wl[17124], wl[17125], wl[17126], wl[17127], wl[17128], wl[17129], wl[17130], wl[17131], wl[17132], wl[17133], wl[17134], wl[17135], wl[17136], wl[17137], wl[17138], wl[17139], wl[17140], wl[17141], wl[17142], wl[17143], wl[17144], wl[17145], wl[17146], wl[17147], wl[17148], wl[17149], wl[17150], wl[17151], wl[17152], wl[17153], wl[17154], wl[17155], wl[17156], wl[17157], wl[17158], wl[17159], wl[17160], wl[17161], wl[17162], wl[17163], wl[17164], wl[17165], wl[17166], wl[17167], wl[17168], wl[17169], wl[17170], wl[17171], wl[17172], wl[17173], wl[17174], wl[17175], wl[17176], wl[17177], wl[17178], wl[17179], wl[17180], wl[17181], wl[17182], wl[17183], wl[17184], wl[17185], wl[17186], wl[17187], wl[17188], wl[17189], wl[17190], wl[17191], wl[17192], wl[17193], wl[17194], wl[17195], wl[17196], wl[17197], wl[17198], wl[17199], wl[17200], wl[17201], wl[17202], wl[17203], wl[17204], wl[17205], wl[17206], wl[17207], wl[17208], wl[17209], wl[17210], wl[17211], wl[17212], wl[17213], wl[17214], wl[17215], wl[17216], wl[17217], wl[17218], wl[17219], wl[17220], wl[17221], wl[17222], wl[17223], wl[17224], wl[17225], wl[17226], wl[17227], wl[17228], wl[17229], wl[17230], wl[17231], wl[17232], wl[17233], wl[17234], wl[17235], wl[17236], wl[17237], wl[17238], wl[17239], wl[17240], wl[17241], wl[17242], wl[17243], wl[17244], wl[17245], wl[17246], wl[17247], wl[17248], wl[17249], wl[17250], wl[17251], wl[17252], wl[17253], wl[17254], wl[17255], wl[17256], wl[17257], wl[17258], wl[17259], wl[17260], wl[17261], wl[17262], wl[17263], wl[17264], wl[17265], wl[17266], wl[17267], wl[17268], wl[17269], wl[17270], wl[17271], wl[17272], wl[17273], wl[17274], wl[17275], wl[17276], wl[17277], wl[17278], wl[17279], wl[17280], wl[17281], wl[17282], wl[17283], wl[17284], wl[17285], wl[17286], wl[17287], wl[17288], wl[17289], wl[17290], wl[17291], wl[17292], wl[17293], wl[17294], wl[17295], wl[17296], wl[17297], wl[17298], wl[17299], wl[17300], wl[17301], wl[17302], wl[17303], wl[17304], wl[17305], wl[17306], wl[17307], wl[17308], wl[17309], wl[17310], wl[17311], wl[17312], wl[17313], wl[17314], wl[17315], wl[17316], wl[17317], wl[17318], wl[17319], wl[17320], wl[17321], wl[17322], wl[17323], wl[17324], wl[17325], wl[17326], wl[17327], wl[17328], wl[17329], wl[17330], wl[17331], wl[17332], wl[17333], wl[17334], wl[17335], wl[17336], wl[17337], wl[17338], wl[17339], wl[17340], wl[17341], wl[17342], wl[17343], wl[17344], wl[17345], wl[17346], wl[17347], wl[17348], wl[17349], wl[17350], wl[17351], wl[17352], wl[17353], wl[17354], wl[17355], wl[17356], wl[17357], wl[17358], wl[17359], wl[17360], wl[17361], wl[17362], wl[17363], wl[17364], wl[17365], wl[17366], wl[17367], wl[17368], wl[17369], wl[17370], wl[17371], wl[17372], wl[17373], wl[17374], wl[17375], wl[17376], wl[17377], wl[17378], wl[17379], wl[17380], wl[17381], wl[17382], wl[17383], wl[17384], wl[17385], wl[17386], wl[17387], wl[17388], wl[17389], wl[17390], wl[17391], wl[17392], wl[17393], wl[17394], wl[17395], wl[17396], wl[17397], wl[17398], wl[17399], wl[17400], wl[17401], wl[17402], wl[17403], wl[17404], wl[17405], wl[17406], wl[17407], wl[17408], wl[17409], wl[17410], wl[17411], wl[17412], wl[17413], wl[17414], wl[17415], wl[17416], wl[17417], wl[17418], wl[17419], wl[17420], wl[17421], wl[17422], wl[17423], wl[17424], wl[17425], wl[17426], wl[17427], wl[17428], wl[17429], wl[17430], wl[17431], wl[17432], wl[17433], wl[17434], wl[17435], wl[17436], wl[17437], wl[17438], wl[17439], wl[17440], wl[17441], wl[17442], wl[17443], wl[17444], wl[17445], wl[17446], wl[17447], wl[17448], wl[17449], wl[17450], wl[17451], wl[17452], wl[17453], wl[17454], wl[17455], wl[17456], wl[17457], wl[17458], wl[17459], wl[17460], wl[17461], wl[17462], wl[17463], wl[17464], wl[17465], wl[17466], wl[17467], wl[17468], wl[17469], wl[17470], wl[17471], wl[17472], wl[17473], wl[17474], wl[17475], wl[17476], wl[17477], wl[17478], wl[17479], wl[17480], wl[17481], wl[17482], wl[17483], wl[17484], wl[17485], wl[17486], wl[17487], wl[17488], wl[17489], wl[17490], wl[17491], wl[17492], wl[17493], wl[17494], wl[17495], wl[17496], wl[17497], wl[17498], wl[17499], wl[17500], wl[17501], wl[17502], wl[17503], wl[17504], wl[17505], wl[17506], wl[17507], wl[17508], wl[17509], wl[17510], wl[17511], wl[17512], wl[17513], wl[17514], wl[17515], wl[17516], wl[17517], wl[17518], wl[17519], wl[17520], wl[17521], wl[17522], wl[17523], wl[17524], wl[17525], wl[17526], wl[17527], wl[17528], wl[17529], wl[17530], wl[17531], wl[17532], wl[17533], wl[17534], wl[17535], wl[17536], wl[17537], wl[17538], wl[17539], wl[17540], wl[17541], wl[17542], wl[17543], wl[17544], wl[17545], wl[17546], wl[17547], wl[17548], wl[17549], wl[17550], wl[17551], wl[17552], wl[17553], wl[17554], wl[17555], wl[17556], wl[17557], wl[17558], wl[17559], wl[17560], wl[17561], wl[17562], wl[17563], wl[17564], wl[17565], wl[17566], wl[17567], wl[17568], wl[17569], wl[17570], wl[17571], wl[17572], wl[17573], wl[17574], wl[17575], wl[17576], wl[17577], wl[17578], wl[17579], wl[17580], wl[17581], wl[17582], wl[17583], wl[17584], wl[17585], wl[17586], wl[17587], wl[17588], wl[17589], wl[17590], wl[17591], wl[17592], wl[17593], wl[17594], wl[17595], wl[17596], wl[17597], wl[17598], wl[17599], wl[17600], wl[17601], wl[17602], wl[17603], wl[17604], wl[17605], wl[17606], wl[17607], wl[17608], wl[17609], wl[17610], wl[17611], wl[17612], wl[17613], wl[17614], wl[17615], wl[17616], wl[17617], wl[17618], wl[17619], wl[17620], wl[17621], wl[17622], wl[17623], wl[17624], wl[17625], wl[17626], wl[17627], wl[17628], wl[17629], wl[17630], wl[17631], wl[17632], wl[17633], wl[17634], wl[17635], wl[17636], wl[17637], wl[17638], wl[17639], wl[17640], wl[17641], wl[17642], wl[17643], wl[17644], wl[17645], wl[17646], wl[17647], wl[17648], wl[17649], wl[17650], wl[17651], wl[17652], wl[17653], wl[17654], wl[17655], wl[17656], wl[17657], wl[17658], wl[17659], wl[17660], wl[17661], wl[17662], wl[17663], wl[17664], wl[17665], wl[17666], wl[17667], wl[17668], wl[17669], wl[17670], wl[17671], wl[17672], wl[17673], wl[17674], wl[17675], wl[17676], wl[17677], wl[17678], wl[17679], wl[17680], wl[17681], wl[17682], wl[17683], wl[17684], wl[17685], wl[17686], wl[17687], wl[17688], wl[17689], wl[17690], wl[17691], wl[17692], wl[17693], wl[17694], wl[17695], wl[17696], wl[17697], wl[17698], wl[17699], wl[17700], wl[17701], wl[17702], wl[17703], wl[17704], wl[17705], wl[17706], wl[17707], wl[17708], wl[17709], wl[17710], wl[17711], wl[17712], wl[17713], wl[17714], wl[17715], wl[17716], wl[17717], wl[17718], wl[17719], wl[17720], wl[17721], wl[17722], wl[17723], wl[17724], wl[17725], wl[17726], wl[17727], wl[216], wl[217], wl[218], wl[219], wl[220], wl[221], wl[222], wl[223], wl[144], wl[145], wl[146], wl[147], wl[148], wl[149], wl[150], wl[151], wl[152], wl[153], wl[154], wl[155], wl[156], wl[157], wl[158], wl[159], wl[160], wl[161], wl[162], wl[163], wl[164], wl[165], wl[166], wl[167], wl[168], wl[169], wl[170], wl[171], wl[172], wl[173], wl[174], wl[175], wl[176], wl[177], wl[178], wl[179], wl[180], wl[181], wl[182], wl[183], wl[184], wl[185], wl[186], wl[187], wl[188], wl[189], wl[190], wl[191], wl[192], wl[193], wl[194], wl[195], wl[196], wl[197], wl[198], wl[199], wl[200], wl[201], wl[202], wl[203], wl[204], wl[205], wl[206], wl[207], wl[208], wl[209], wl[210], wl[211], wl[212], wl[213], wl[214], wl[215], wl[56], wl[57], wl[58], wl[59], wl[60], wl[61], wl[62], wl[63], wl[16636], wl[16637], wl[16638], wl[16639], wl[16640], wl[16641], wl[16642], wl[16643], wl[16644], wl[16645], wl[16646], wl[16647], wl[16648], wl[16649], wl[16650], wl[16651], wl[16652], wl[16653], wl[16654], wl[16655], wl[16656], wl[16657], wl[16658], wl[16659], wl[16660], wl[16661], wl[16662], wl[16663], wl[16664], wl[16665], wl[16666], wl[16667], wl[16668], wl[16669], wl[16670], wl[16671], wl[16672], wl[16673], wl[16674], wl[16675], wl[16676], wl[16677], wl[16678], wl[16679], wl[16680], wl[16681], wl[16682], wl[16683], wl[16684], wl[16685], wl[16686], wl[16687], wl[16688], wl[16689], wl[16690], wl[16691], wl[16692], wl[16693], wl[16694], wl[16695], wl[16696], wl[16697], wl[16698], wl[16699], wl[16700], wl[16701], wl[16702], wl[16703], wl[16704], wl[16705], wl[16706], wl[16707], wl[64], wl[65], wl[66], wl[67], wl[68], wl[69], wl[70], wl[71], wl[72], wl[73], wl[74], wl[75], wl[76], wl[77], wl[78], wl[79], wl[80], wl[81], wl[82], wl[83], wl[84], wl[85], wl[86], wl[87], wl[88], wl[89], wl[90], wl[91], wl[92], wl[93], wl[94], wl[95], wl[96], wl[97], wl[98], wl[99], wl[100], wl[101], wl[102], wl[103], wl[104], wl[105], wl[106], wl[107], wl[108], wl[109], wl[110], wl[111], wl[112], wl[113], wl[114], wl[115], wl[116], wl[117], wl[118], wl[119], wl[120], wl[121], wl[122], wl[123], wl[124], wl[125], wl[126], wl[127], wl[128], wl[129], wl[130], wl[131], wl[132], wl[133], wl[134], wl[135], wl[136], wl[137], wl[138], wl[139], wl[140], wl[141], wl[142], wl[143]})
    );
    bottom_left_tile tile_1__1_
    (
        .chany_top_in(cby_0__1__0_chany_bottom_out),
        .chanx_right_in(cbx_1__0__0_chanx_left_out),
        .chany_top_out(sb_0__0__0_chany_top_out),
        .chanx_right_out(sb_0__0__0_chanx_right_out),
        .grid_top_r_in(sb_0__0__grid_top_r_in),
        .grid_top_l_inpad(grid_io_left_0__1__io_right_in),
        .grid_right_t_in(sb_0__0__grid_right_t_in),
        .grid_right_b_inpad(grid_io_bottom_1__0__io_top_in),
        .bl(bl[1258:1337]),
        .wl(wl[1258:1337])
    );
    bottom_right_tile tile_5__1_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[64:71]),
        .io_top_in(grid_io_bottom_4__0__io_top_in),
        .chanx_left_in(sb_1__0__2_chanx_right_out),
        .chanx_left_out(cbx_1__0__3_chanx_left_out),
        .grid_top_out(grid_clb_4__1__grid_bottom_in),
        .chany_top_in(cby_4__1__0_chany_bottom_out),
        .chany_top_out(sb_4__0__0_chany_top_out),
        .grid_top_r_inpad(grid_io_right_5__1__io_left_in),
        .grid_top_l_in(sb_4__0__grid_top_l_in),
        .grid_left_t_in(sb_3__0__grid_right_t_in),
        .bl({bl[24], bl[25], bl[26], bl[27], bl[28], bl[29], bl[30], bl[31], bl[5248], bl[5249], bl[5250], bl[5251], bl[5252], bl[5253], bl[5254], bl[5255], bl[5256], bl[5257], bl[5258], bl[5259], bl[5260], bl[5261], bl[5262], bl[5263], bl[5264], bl[5265], bl[5266], bl[5267], bl[5268], bl[5269], bl[5270], bl[5271], bl[5272], bl[5273], bl[5274], bl[5275], bl[5276], bl[5277], bl[5278], bl[5279], bl[5280], bl[5281], bl[5282], bl[5283], bl[5284], bl[5285], bl[5286], bl[5287], bl[5288], bl[5289], bl[5290], bl[5291], bl[5292], bl[5293], bl[5294], bl[5295], bl[5296], bl[5297], bl[5298], bl[5299], bl[5300], bl[5301], bl[5302], bl[5303], bl[5304], bl[5305], bl[5306], bl[5307], bl[5308], bl[5309], bl[5310], bl[5311], bl[5312], bl[5313], bl[5314], bl[5315], bl[5316], bl[5317], bl[5318], bl[5319], bl[5168], bl[5169], bl[5170], bl[5171], bl[5172], bl[5173], bl[5174], bl[5175], bl[5176], bl[5177], bl[5178], bl[5179], bl[5180], bl[5181], bl[5182], bl[5183], bl[5184], bl[5185], bl[5186], bl[5187], bl[5188], bl[5189], bl[5190], bl[5191], bl[5192], bl[5193], bl[5194], bl[5195], bl[5196], bl[5197], bl[5198], bl[5199], bl[5200], bl[5201], bl[5202], bl[5203], bl[5204], bl[5205], bl[5206], bl[5207], bl[5208], bl[5209], bl[5210], bl[5211], bl[5212], bl[5213], bl[5214], bl[5215], bl[5216], bl[5217], bl[5218], bl[5219], bl[5220], bl[5221], bl[5222], bl[5223], bl[5224], bl[5225], bl[5226], bl[5227], bl[5228], bl[5229], bl[5230], bl[5231], bl[5232], bl[5233], bl[5234], bl[5235], bl[5236], bl[5237], bl[5238], bl[5239], bl[5240], bl[5241], bl[5242], bl[5243], bl[5244], bl[5245], bl[5246], bl[5247]}),
        .wl({wl[24], wl[25], wl[26], wl[27], wl[28], wl[29], wl[30], wl[31], wl[5248], wl[5249], wl[5250], wl[5251], wl[5252], wl[5253], wl[5254], wl[5255], wl[5256], wl[5257], wl[5258], wl[5259], wl[5260], wl[5261], wl[5262], wl[5263], wl[5264], wl[5265], wl[5266], wl[5267], wl[5268], wl[5269], wl[5270], wl[5271], wl[5272], wl[5273], wl[5274], wl[5275], wl[5276], wl[5277], wl[5278], wl[5279], wl[5280], wl[5281], wl[5282], wl[5283], wl[5284], wl[5285], wl[5286], wl[5287], wl[5288], wl[5289], wl[5290], wl[5291], wl[5292], wl[5293], wl[5294], wl[5295], wl[5296], wl[5297], wl[5298], wl[5299], wl[5300], wl[5301], wl[5302], wl[5303], wl[5304], wl[5305], wl[5306], wl[5307], wl[5308], wl[5309], wl[5310], wl[5311], wl[5312], wl[5313], wl[5314], wl[5315], wl[5316], wl[5317], wl[5318], wl[5319], wl[5168], wl[5169], wl[5170], wl[5171], wl[5172], wl[5173], wl[5174], wl[5175], wl[5176], wl[5177], wl[5178], wl[5179], wl[5180], wl[5181], wl[5182], wl[5183], wl[5184], wl[5185], wl[5186], wl[5187], wl[5188], wl[5189], wl[5190], wl[5191], wl[5192], wl[5193], wl[5194], wl[5195], wl[5196], wl[5197], wl[5198], wl[5199], wl[5200], wl[5201], wl[5202], wl[5203], wl[5204], wl[5205], wl[5206], wl[5207], wl[5208], wl[5209], wl[5210], wl[5211], wl[5212], wl[5213], wl[5214], wl[5215], wl[5216], wl[5217], wl[5218], wl[5219], wl[5220], wl[5221], wl[5222], wl[5223], wl[5224], wl[5225], wl[5226], wl[5227], wl[5228], wl[5229], wl[5230], wl[5231], wl[5232], wl[5233], wl[5234], wl[5235], wl[5236], wl[5237], wl[5238], wl[5239], wl[5240], wl[5241], wl[5242], wl[5243], wl[5244], wl[5245], wl[5246], wl[5247]})
    );
    left_tile tile_1__2_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[96:103]),
        .io_right_in(grid_io_left_0__1__io_right_in),
        .chany_bottom_in(sb_0__0__0_chany_top_out),
        .chany_bottom_out(cby_0__1__0_chany_bottom_out),
        .grid_right_out(grid_clb_1__1__grid_left_in),
        .chany_top_in_0(cby_0__1__1_chany_bottom_out),
        .chanx_right_in(cbx_1__1__0_chanx_left_out),
        .chany_top_out_0(sb_0__1__0_chany_top_out),
        .chanx_right_out(sb_0__1__0_chanx_right_out),
        .grid_top_r_in(sb_0__1__grid_top_r_in),
        .grid_top_l_inpad(grid_io_left_0__2__io_right_in),
        .grid_right_t_in(sb_0__1__grid_right_t_in),
        .grid_right_b_in(sb_0__1__grid_right_b_in),
        .grid_bottom_r_in(sb_0__0__grid_top_r_in),
        .bl({bl[1410], bl[1411], bl[1412], bl[1413], bl[1414], bl[1415], bl[1416], bl[1417], bl[1338], bl[1339], bl[1340], bl[1341], bl[1342], bl[1343], bl[1344], bl[1345], bl[1346], bl[1347], bl[1348], bl[1349], bl[1350], bl[1351], bl[1352], bl[1353], bl[1354], bl[1355], bl[1356], bl[1357], bl[1358], bl[1359], bl[1360], bl[1361], bl[1362], bl[1363], bl[1364], bl[1365], bl[1366], bl[1367], bl[1368], bl[1369], bl[1370], bl[1371], bl[1372], bl[1373], bl[1374], bl[1375], bl[1376], bl[1377], bl[1378], bl[1379], bl[1380], bl[1381], bl[1382], bl[1383], bl[1384], bl[1385], bl[1386], bl[1387], bl[1388], bl[1389], bl[1390], bl[1391], bl[1392], bl[1393], bl[1394], bl[1395], bl[1396], bl[1397], bl[1398], bl[1399], bl[1400], bl[1401], bl[1402], bl[1403], bl[1404], bl[1405], bl[1406], bl[1407], bl[1408], bl[1409], bl[1100], bl[1101], bl[1102], bl[1103], bl[1104], bl[1105], bl[1106], bl[1107], bl[1108], bl[1109], bl[1110], bl[1111], bl[1112], bl[1113], bl[1114], bl[1115], bl[1116], bl[1117], bl[1118], bl[1119], bl[1120], bl[1121], bl[1122], bl[1123], bl[1124], bl[1125], bl[1126], bl[1127], bl[1128], bl[1129], bl[1130], bl[1131], bl[1132], bl[1133], bl[1134], bl[1135], bl[1136], bl[1137], bl[1138], bl[1139], bl[1140], bl[1141], bl[1142], bl[1143], bl[1144], bl[1145], bl[1146], bl[1147], bl[1148], bl[1149], bl[1150], bl[1151], bl[1152], bl[1153], bl[1154], bl[1155], bl[1156], bl[1157], bl[1158], bl[1159], bl[1160], bl[1161], bl[1162], bl[1163], bl[1164], bl[1165], bl[1166], bl[1167], bl[1168], bl[1169], bl[1170], bl[1171], bl[1172], bl[1173], bl[1174], bl[1175], bl[1176], bl[1177]}),
        .wl({wl[1410], wl[1411], wl[1412], wl[1413], wl[1414], wl[1415], wl[1416], wl[1417], wl[1338], wl[1339], wl[1340], wl[1341], wl[1342], wl[1343], wl[1344], wl[1345], wl[1346], wl[1347], wl[1348], wl[1349], wl[1350], wl[1351], wl[1352], wl[1353], wl[1354], wl[1355], wl[1356], wl[1357], wl[1358], wl[1359], wl[1360], wl[1361], wl[1362], wl[1363], wl[1364], wl[1365], wl[1366], wl[1367], wl[1368], wl[1369], wl[1370], wl[1371], wl[1372], wl[1373], wl[1374], wl[1375], wl[1376], wl[1377], wl[1378], wl[1379], wl[1380], wl[1381], wl[1382], wl[1383], wl[1384], wl[1385], wl[1386], wl[1387], wl[1388], wl[1389], wl[1390], wl[1391], wl[1392], wl[1393], wl[1394], wl[1395], wl[1396], wl[1397], wl[1398], wl[1399], wl[1400], wl[1401], wl[1402], wl[1403], wl[1404], wl[1405], wl[1406], wl[1407], wl[1408], wl[1409], wl[1100], wl[1101], wl[1102], wl[1103], wl[1104], wl[1105], wl[1106], wl[1107], wl[1108], wl[1109], wl[1110], wl[1111], wl[1112], wl[1113], wl[1114], wl[1115], wl[1116], wl[1117], wl[1118], wl[1119], wl[1120], wl[1121], wl[1122], wl[1123], wl[1124], wl[1125], wl[1126], wl[1127], wl[1128], wl[1129], wl[1130], wl[1131], wl[1132], wl[1133], wl[1134], wl[1135], wl[1136], wl[1137], wl[1138], wl[1139], wl[1140], wl[1141], wl[1142], wl[1143], wl[1144], wl[1145], wl[1146], wl[1147], wl[1148], wl[1149], wl[1150], wl[1151], wl[1152], wl[1153], wl[1154], wl[1155], wl[1156], wl[1157], wl[1158], wl[1159], wl[1160], wl[1161], wl[1162], wl[1163], wl[1164], wl[1165], wl[1166], wl[1167], wl[1168], wl[1169], wl[1170], wl[1171], wl[1172], wl[1173], wl[1174], wl[1175], wl[1176], wl[1177]})
    );
    left_tile tile_1__3_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[104:111]),
        .io_right_in(grid_io_left_0__2__io_right_in),
        .chany_bottom_in(sb_0__1__0_chany_top_out),
        .chany_bottom_out(cby_0__1__1_chany_bottom_out),
        .grid_right_out(grid_clb_1__2__grid_left_in),
        .chany_top_in_0(cby_0__1__2_chany_bottom_out),
        .chanx_right_in(cbx_1__1__1_chanx_left_out),
        .chany_top_out_0(sb_0__1__1_chany_top_out),
        .chanx_right_out(sb_0__1__1_chanx_right_out),
        .grid_top_r_in(sb_0__2__grid_top_r_in),
        .grid_top_l_inpad(grid_io_left_0__3__io_right_in),
        .grid_right_t_in(sb_0__2__grid_right_t_in),
        .grid_right_b_in(sb_0__2__grid_right_b_in),
        .grid_bottom_r_in(sb_0__1__grid_top_r_in),
        .bl({bl[1250], bl[1251], bl[1252], bl[1253], bl[1254], bl[1255], bl[1256], bl[1257], bl[1178], bl[1179], bl[1180], bl[1181], bl[1182], bl[1183], bl[1184], bl[1185], bl[1186], bl[1187], bl[1188], bl[1189], bl[1190], bl[1191], bl[1192], bl[1193], bl[1194], bl[1195], bl[1196], bl[1197], bl[1198], bl[1199], bl[1200], bl[1201], bl[1202], bl[1203], bl[1204], bl[1205], bl[1206], bl[1207], bl[1208], bl[1209], bl[1210], bl[1211], bl[1212], bl[1213], bl[1214], bl[1215], bl[1216], bl[1217], bl[1218], bl[1219], bl[1220], bl[1221], bl[1222], bl[1223], bl[1224], bl[1225], bl[1226], bl[1227], bl[1228], bl[1229], bl[1230], bl[1231], bl[1232], bl[1233], bl[1234], bl[1235], bl[1236], bl[1237], bl[1238], bl[1239], bl[1240], bl[1241], bl[1242], bl[1243], bl[1244], bl[1245], bl[1246], bl[1247], bl[1248], bl[1249], bl[942], bl[943], bl[944], bl[945], bl[946], bl[947], bl[948], bl[949], bl[950], bl[951], bl[952], bl[953], bl[954], bl[955], bl[956], bl[957], bl[958], bl[959], bl[960], bl[961], bl[962], bl[963], bl[964], bl[965], bl[966], bl[967], bl[968], bl[969], bl[970], bl[971], bl[972], bl[973], bl[974], bl[975], bl[976], bl[977], bl[978], bl[979], bl[980], bl[981], bl[982], bl[983], bl[984], bl[985], bl[986], bl[987], bl[988], bl[989], bl[990], bl[991], bl[992], bl[993], bl[994], bl[995], bl[996], bl[997], bl[998], bl[999], bl[1000], bl[1001], bl[1002], bl[1003], bl[1004], bl[1005], bl[1006], bl[1007], bl[1008], bl[1009], bl[1010], bl[1011], bl[1012], bl[1013], bl[1014], bl[1015], bl[1016], bl[1017], bl[1018], bl[1019]}),
        .wl({wl[1250], wl[1251], wl[1252], wl[1253], wl[1254], wl[1255], wl[1256], wl[1257], wl[1178], wl[1179], wl[1180], wl[1181], wl[1182], wl[1183], wl[1184], wl[1185], wl[1186], wl[1187], wl[1188], wl[1189], wl[1190], wl[1191], wl[1192], wl[1193], wl[1194], wl[1195], wl[1196], wl[1197], wl[1198], wl[1199], wl[1200], wl[1201], wl[1202], wl[1203], wl[1204], wl[1205], wl[1206], wl[1207], wl[1208], wl[1209], wl[1210], wl[1211], wl[1212], wl[1213], wl[1214], wl[1215], wl[1216], wl[1217], wl[1218], wl[1219], wl[1220], wl[1221], wl[1222], wl[1223], wl[1224], wl[1225], wl[1226], wl[1227], wl[1228], wl[1229], wl[1230], wl[1231], wl[1232], wl[1233], wl[1234], wl[1235], wl[1236], wl[1237], wl[1238], wl[1239], wl[1240], wl[1241], wl[1242], wl[1243], wl[1244], wl[1245], wl[1246], wl[1247], wl[1248], wl[1249], wl[942], wl[943], wl[944], wl[945], wl[946], wl[947], wl[948], wl[949], wl[950], wl[951], wl[952], wl[953], wl[954], wl[955], wl[956], wl[957], wl[958], wl[959], wl[960], wl[961], wl[962], wl[963], wl[964], wl[965], wl[966], wl[967], wl[968], wl[969], wl[970], wl[971], wl[972], wl[973], wl[974], wl[975], wl[976], wl[977], wl[978], wl[979], wl[980], wl[981], wl[982], wl[983], wl[984], wl[985], wl[986], wl[987], wl[988], wl[989], wl[990], wl[991], wl[992], wl[993], wl[994], wl[995], wl[996], wl[997], wl[998], wl[999], wl[1000], wl[1001], wl[1002], wl[1003], wl[1004], wl[1005], wl[1006], wl[1007], wl[1008], wl[1009], wl[1010], wl[1011], wl[1012], wl[1013], wl[1014], wl[1015], wl[1016], wl[1017], wl[1018], wl[1019]})
    );
    left_tile tile_1__4_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[112:119]),
        .io_right_in(grid_io_left_0__3__io_right_in),
        .chany_bottom_in(sb_0__1__1_chany_top_out),
        .chany_bottom_out(cby_0__1__2_chany_bottom_out),
        .grid_right_out(grid_clb_1__3__grid_left_in),
        .chany_top_in_0(cby_0__1__3_chany_bottom_out),
        .chanx_right_in(cbx_1__1__2_chanx_left_out),
        .chany_top_out_0(sb_0__1__2_chany_top_out),
        .chanx_right_out(sb_0__1__2_chanx_right_out),
        .grid_top_r_in(sb_0__3__grid_top_r_in),
        .grid_top_l_inpad(grid_io_left_0__4__io_right_in),
        .grid_right_t_in(sb_0__3__grid_right_t_in),
        .grid_right_b_in(sb_0__3__grid_right_b_in),
        .grid_bottom_r_in(sb_0__2__grid_top_r_in),
        .bl({bl[1092], bl[1093], bl[1094], bl[1095], bl[1096], bl[1097], bl[1098], bl[1099], bl[1020], bl[1021], bl[1022], bl[1023], bl[1024], bl[1025], bl[1026], bl[1027], bl[1028], bl[1029], bl[1030], bl[1031], bl[1032], bl[1033], bl[1034], bl[1035], bl[1036], bl[1037], bl[1038], bl[1039], bl[1040], bl[1041], bl[1042], bl[1043], bl[1044], bl[1045], bl[1046], bl[1047], bl[1048], bl[1049], bl[1050], bl[1051], bl[1052], bl[1053], bl[1054], bl[1055], bl[1056], bl[1057], bl[1058], bl[1059], bl[1060], bl[1061], bl[1062], bl[1063], bl[1064], bl[1065], bl[1066], bl[1067], bl[1068], bl[1069], bl[1070], bl[1071], bl[1072], bl[1073], bl[1074], bl[1075], bl[1076], bl[1077], bl[1078], bl[1079], bl[1080], bl[1081], bl[1082], bl[1083], bl[1084], bl[1085], bl[1086], bl[1087], bl[1088], bl[1089], bl[1090], bl[1091], bl[784], bl[785], bl[786], bl[787], bl[788], bl[789], bl[790], bl[791], bl[792], bl[793], bl[794], bl[795], bl[796], bl[797], bl[798], bl[799], bl[800], bl[801], bl[802], bl[803], bl[804], bl[805], bl[806], bl[807], bl[808], bl[809], bl[810], bl[811], bl[812], bl[813], bl[814], bl[815], bl[816], bl[817], bl[818], bl[819], bl[820], bl[821], bl[822], bl[823], bl[824], bl[825], bl[826], bl[827], bl[828], bl[829], bl[830], bl[831], bl[832], bl[833], bl[834], bl[835], bl[836], bl[837], bl[838], bl[839], bl[840], bl[841], bl[842], bl[843], bl[844], bl[845], bl[846], bl[847], bl[848], bl[849], bl[850], bl[851], bl[852], bl[853], bl[854], bl[855], bl[856], bl[857], bl[858], bl[859], bl[860], bl[861]}),
        .wl({wl[1092], wl[1093], wl[1094], wl[1095], wl[1096], wl[1097], wl[1098], wl[1099], wl[1020], wl[1021], wl[1022], wl[1023], wl[1024], wl[1025], wl[1026], wl[1027], wl[1028], wl[1029], wl[1030], wl[1031], wl[1032], wl[1033], wl[1034], wl[1035], wl[1036], wl[1037], wl[1038], wl[1039], wl[1040], wl[1041], wl[1042], wl[1043], wl[1044], wl[1045], wl[1046], wl[1047], wl[1048], wl[1049], wl[1050], wl[1051], wl[1052], wl[1053], wl[1054], wl[1055], wl[1056], wl[1057], wl[1058], wl[1059], wl[1060], wl[1061], wl[1062], wl[1063], wl[1064], wl[1065], wl[1066], wl[1067], wl[1068], wl[1069], wl[1070], wl[1071], wl[1072], wl[1073], wl[1074], wl[1075], wl[1076], wl[1077], wl[1078], wl[1079], wl[1080], wl[1081], wl[1082], wl[1083], wl[1084], wl[1085], wl[1086], wl[1087], wl[1088], wl[1089], wl[1090], wl[1091], wl[784], wl[785], wl[786], wl[787], wl[788], wl[789], wl[790], wl[791], wl[792], wl[793], wl[794], wl[795], wl[796], wl[797], wl[798], wl[799], wl[800], wl[801], wl[802], wl[803], wl[804], wl[805], wl[806], wl[807], wl[808], wl[809], wl[810], wl[811], wl[812], wl[813], wl[814], wl[815], wl[816], wl[817], wl[818], wl[819], wl[820], wl[821], wl[822], wl[823], wl[824], wl[825], wl[826], wl[827], wl[828], wl[829], wl[830], wl[831], wl[832], wl[833], wl[834], wl[835], wl[836], wl[837], wl[838], wl[839], wl[840], wl[841], wl[842], wl[843], wl[844], wl[845], wl[846], wl[847], wl[848], wl[849], wl[850], wl[851], wl[852], wl[853], wl[854], wl[855], wl[856], wl[857], wl[858], wl[859], wl[860], wl[861]})
    );
    bottom_tile tile_2__1_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[88:95]),
        .io_top_in(grid_io_bottom_1__0__io_top_in),
        .chanx_left_in(sb_0__0__0_chanx_right_out),
        .chanx_left_out(cbx_1__0__0_chanx_left_out),
        .grid_top_out(grid_clb_1__1__grid_bottom_in),
        .chany_top_in(cby_1__1__0_chany_bottom_out),
        .chanx_right_in_0(cbx_1__0__1_chanx_left_out),
        .chany_top_out(sb_1__0__0_chany_top_out),
        .chanx_right_out_0(sb_1__0__0_chanx_right_out),
        .grid_top_r_in(sb_1__0__grid_top_r_in),
        .grid_top_l_in(sb_1__0__grid_top_l_in),
        .grid_right_t_in(sb_1__0__grid_right_t_in),
        .grid_right_b_inpad(grid_io_bottom_2__0__io_top_in),
        .grid_left_t_in(sb_0__0__grid_right_t_in),
        .bl({bl[0], bl[1], bl[2], bl[3], bl[4], bl[5], bl[6], bl[7], bl[1496], bl[1497], bl[1498], bl[1499], bl[1500], bl[1501], bl[1502], bl[1503], bl[1504], bl[1505], bl[1506], bl[1507], bl[1508], bl[1509], bl[1510], bl[1511], bl[1512], bl[1513], bl[1514], bl[1515], bl[1516], bl[1517], bl[1518], bl[1519], bl[1520], bl[1521], bl[1522], bl[1523], bl[1524], bl[1525], bl[1526], bl[1527], bl[1528], bl[1529], bl[1530], bl[1531], bl[1532], bl[1533], bl[1534], bl[1535], bl[1536], bl[1537], bl[1538], bl[1539], bl[1540], bl[1541], bl[1542], bl[1543], bl[1544], bl[1545], bl[1546], bl[1547], bl[1548], bl[1549], bl[1550], bl[1551], bl[1552], bl[1553], bl[1554], bl[1555], bl[1556], bl[1557], bl[1558], bl[1559], bl[1560], bl[1561], bl[1562], bl[1563], bl[1564], bl[1565], bl[1566], bl[1567], bl[1418], bl[1419], bl[1420], bl[1421], bl[1422], bl[1423], bl[1424], bl[1425], bl[1426], bl[1427], bl[1428], bl[1429], bl[1430], bl[1431], bl[1432], bl[1433], bl[1434], bl[1435], bl[1436], bl[1437], bl[1438], bl[1439], bl[1440], bl[1441], bl[1442], bl[1443], bl[1444], bl[1445], bl[1446], bl[1447], bl[1448], bl[1449], bl[1450], bl[1451], bl[1452], bl[1453], bl[1454], bl[1455], bl[1456], bl[1457], bl[1458], bl[1459], bl[1460], bl[1461], bl[1462], bl[1463], bl[1464], bl[1465], bl[1466], bl[1467], bl[1468], bl[1469], bl[1470], bl[1471], bl[1472], bl[1473], bl[1474], bl[1475], bl[1476], bl[1477], bl[1478], bl[1479], bl[1480], bl[1481], bl[1482], bl[1483], bl[1484], bl[1485], bl[1486], bl[1487], bl[1488], bl[1489], bl[1490], bl[1491], bl[1492], bl[1493], bl[1494], bl[1495]}),
        .wl({wl[0], wl[1], wl[2], wl[3], wl[4], wl[5], wl[6], wl[7], wl[1496], wl[1497], wl[1498], wl[1499], wl[1500], wl[1501], wl[1502], wl[1503], wl[1504], wl[1505], wl[1506], wl[1507], wl[1508], wl[1509], wl[1510], wl[1511], wl[1512], wl[1513], wl[1514], wl[1515], wl[1516], wl[1517], wl[1518], wl[1519], wl[1520], wl[1521], wl[1522], wl[1523], wl[1524], wl[1525], wl[1526], wl[1527], wl[1528], wl[1529], wl[1530], wl[1531], wl[1532], wl[1533], wl[1534], wl[1535], wl[1536], wl[1537], wl[1538], wl[1539], wl[1540], wl[1541], wl[1542], wl[1543], wl[1544], wl[1545], wl[1546], wl[1547], wl[1548], wl[1549], wl[1550], wl[1551], wl[1552], wl[1553], wl[1554], wl[1555], wl[1556], wl[1557], wl[1558], wl[1559], wl[1560], wl[1561], wl[1562], wl[1563], wl[1564], wl[1565], wl[1566], wl[1567], wl[1418], wl[1419], wl[1420], wl[1421], wl[1422], wl[1423], wl[1424], wl[1425], wl[1426], wl[1427], wl[1428], wl[1429], wl[1430], wl[1431], wl[1432], wl[1433], wl[1434], wl[1435], wl[1436], wl[1437], wl[1438], wl[1439], wl[1440], wl[1441], wl[1442], wl[1443], wl[1444], wl[1445], wl[1446], wl[1447], wl[1448], wl[1449], wl[1450], wl[1451], wl[1452], wl[1453], wl[1454], wl[1455], wl[1456], wl[1457], wl[1458], wl[1459], wl[1460], wl[1461], wl[1462], wl[1463], wl[1464], wl[1465], wl[1466], wl[1467], wl[1468], wl[1469], wl[1470], wl[1471], wl[1472], wl[1473], wl[1474], wl[1475], wl[1476], wl[1477], wl[1478], wl[1479], wl[1480], wl[1481], wl[1482], wl[1483], wl[1484], wl[1485], wl[1486], wl[1487], wl[1488], wl[1489], wl[1490], wl[1491], wl[1492], wl[1493], wl[1494], wl[1495]})
    );
    bottom_tile tile_3__1_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[80:87]),
        .io_top_in(grid_io_bottom_2__0__io_top_in),
        .chanx_left_in(sb_1__0__0_chanx_right_out),
        .chanx_left_out(cbx_1__0__1_chanx_left_out),
        .grid_top_out(grid_clb_2__1__grid_bottom_in),
        .chany_top_in(cby_1__1__4_chany_bottom_out),
        .chanx_right_in_0(cbx_1__0__2_chanx_left_out),
        .chany_top_out(sb_1__0__1_chany_top_out),
        .chanx_right_out_0(sb_1__0__1_chanx_right_out),
        .grid_top_r_in(sb_2__0__grid_top_r_in),
        .grid_top_l_in(sb_2__0__grid_top_l_in),
        .grid_right_t_in(sb_2__0__grid_right_t_in),
        .grid_right_b_inpad(grid_io_bottom_3__0__io_top_in),
        .grid_left_t_in(sb_1__0__grid_right_t_in),
        .bl({bl[8], bl[9], bl[10], bl[11], bl[12], bl[13], bl[14], bl[15], bl[2746], bl[2747], bl[2748], bl[2749], bl[2750], bl[2751], bl[2752], bl[2753], bl[2754], bl[2755], bl[2756], bl[2757], bl[2758], bl[2759], bl[2760], bl[2761], bl[2762], bl[2763], bl[2764], bl[2765], bl[2766], bl[2767], bl[2768], bl[2769], bl[2770], bl[2771], bl[2772], bl[2773], bl[2774], bl[2775], bl[2776], bl[2777], bl[2778], bl[2779], bl[2780], bl[2781], bl[2782], bl[2783], bl[2784], bl[2785], bl[2786], bl[2787], bl[2788], bl[2789], bl[2790], bl[2791], bl[2792], bl[2793], bl[2794], bl[2795], bl[2796], bl[2797], bl[2798], bl[2799], bl[2800], bl[2801], bl[2802], bl[2803], bl[2804], bl[2805], bl[2806], bl[2807], bl[2808], bl[2809], bl[2810], bl[2811], bl[2812], bl[2813], bl[2814], bl[2815], bl[2816], bl[2817], bl[2668], bl[2669], bl[2670], bl[2671], bl[2672], bl[2673], bl[2674], bl[2675], bl[2676], bl[2677], bl[2678], bl[2679], bl[2680], bl[2681], bl[2682], bl[2683], bl[2684], bl[2685], bl[2686], bl[2687], bl[2688], bl[2689], bl[2690], bl[2691], bl[2692], bl[2693], bl[2694], bl[2695], bl[2696], bl[2697], bl[2698], bl[2699], bl[2700], bl[2701], bl[2702], bl[2703], bl[2704], bl[2705], bl[2706], bl[2707], bl[2708], bl[2709], bl[2710], bl[2711], bl[2712], bl[2713], bl[2714], bl[2715], bl[2716], bl[2717], bl[2718], bl[2719], bl[2720], bl[2721], bl[2722], bl[2723], bl[2724], bl[2725], bl[2726], bl[2727], bl[2728], bl[2729], bl[2730], bl[2731], bl[2732], bl[2733], bl[2734], bl[2735], bl[2736], bl[2737], bl[2738], bl[2739], bl[2740], bl[2741], bl[2742], bl[2743], bl[2744], bl[2745]}),
        .wl({wl[8], wl[9], wl[10], wl[11], wl[12], wl[13], wl[14], wl[15], wl[2746], wl[2747], wl[2748], wl[2749], wl[2750], wl[2751], wl[2752], wl[2753], wl[2754], wl[2755], wl[2756], wl[2757], wl[2758], wl[2759], wl[2760], wl[2761], wl[2762], wl[2763], wl[2764], wl[2765], wl[2766], wl[2767], wl[2768], wl[2769], wl[2770], wl[2771], wl[2772], wl[2773], wl[2774], wl[2775], wl[2776], wl[2777], wl[2778], wl[2779], wl[2780], wl[2781], wl[2782], wl[2783], wl[2784], wl[2785], wl[2786], wl[2787], wl[2788], wl[2789], wl[2790], wl[2791], wl[2792], wl[2793], wl[2794], wl[2795], wl[2796], wl[2797], wl[2798], wl[2799], wl[2800], wl[2801], wl[2802], wl[2803], wl[2804], wl[2805], wl[2806], wl[2807], wl[2808], wl[2809], wl[2810], wl[2811], wl[2812], wl[2813], wl[2814], wl[2815], wl[2816], wl[2817], wl[2668], wl[2669], wl[2670], wl[2671], wl[2672], wl[2673], wl[2674], wl[2675], wl[2676], wl[2677], wl[2678], wl[2679], wl[2680], wl[2681], wl[2682], wl[2683], wl[2684], wl[2685], wl[2686], wl[2687], wl[2688], wl[2689], wl[2690], wl[2691], wl[2692], wl[2693], wl[2694], wl[2695], wl[2696], wl[2697], wl[2698], wl[2699], wl[2700], wl[2701], wl[2702], wl[2703], wl[2704], wl[2705], wl[2706], wl[2707], wl[2708], wl[2709], wl[2710], wl[2711], wl[2712], wl[2713], wl[2714], wl[2715], wl[2716], wl[2717], wl[2718], wl[2719], wl[2720], wl[2721], wl[2722], wl[2723], wl[2724], wl[2725], wl[2726], wl[2727], wl[2728], wl[2729], wl[2730], wl[2731], wl[2732], wl[2733], wl[2734], wl[2735], wl[2736], wl[2737], wl[2738], wl[2739], wl[2740], wl[2741], wl[2742], wl[2743], wl[2744], wl[2745]})
    );
    bottom_tile tile_4__1_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[72:79]),
        .io_top_in(grid_io_bottom_3__0__io_top_in),
        .chanx_left_in(sb_1__0__1_chanx_right_out),
        .chanx_left_out(cbx_1__0__2_chanx_left_out),
        .grid_top_out(grid_clb_3__1__grid_bottom_in),
        .chany_top_in(cby_1__1__8_chany_bottom_out),
        .chanx_right_in_0(cbx_1__0__3_chanx_left_out),
        .chany_top_out(sb_1__0__2_chany_top_out),
        .chanx_right_out_0(sb_1__0__2_chanx_right_out),
        .grid_top_r_in(sb_3__0__grid_top_r_in),
        .grid_top_l_in(sb_3__0__grid_top_l_in),
        .grid_right_t_in(sb_3__0__grid_right_t_in),
        .grid_right_b_inpad(grid_io_bottom_4__0__io_top_in),
        .grid_left_t_in(sb_2__0__grid_right_t_in),
        .bl({bl[16], bl[17], bl[18], bl[19], bl[20], bl[21], bl[22], bl[23], bl[3996], bl[3997], bl[3998], bl[3999], bl[4000], bl[4001], bl[4002], bl[4003], bl[4004], bl[4005], bl[4006], bl[4007], bl[4008], bl[4009], bl[4010], bl[4011], bl[4012], bl[4013], bl[4014], bl[4015], bl[4016], bl[4017], bl[4018], bl[4019], bl[4020], bl[4021], bl[4022], bl[4023], bl[4024], bl[4025], bl[4026], bl[4027], bl[4028], bl[4029], bl[4030], bl[4031], bl[4032], bl[4033], bl[4034], bl[4035], bl[4036], bl[4037], bl[4038], bl[4039], bl[4040], bl[4041], bl[4042], bl[4043], bl[4044], bl[4045], bl[4046], bl[4047], bl[4048], bl[4049], bl[4050], bl[4051], bl[4052], bl[4053], bl[4054], bl[4055], bl[4056], bl[4057], bl[4058], bl[4059], bl[4060], bl[4061], bl[4062], bl[4063], bl[4064], bl[4065], bl[4066], bl[4067], bl[3918], bl[3919], bl[3920], bl[3921], bl[3922], bl[3923], bl[3924], bl[3925], bl[3926], bl[3927], bl[3928], bl[3929], bl[3930], bl[3931], bl[3932], bl[3933], bl[3934], bl[3935], bl[3936], bl[3937], bl[3938], bl[3939], bl[3940], bl[3941], bl[3942], bl[3943], bl[3944], bl[3945], bl[3946], bl[3947], bl[3948], bl[3949], bl[3950], bl[3951], bl[3952], bl[3953], bl[3954], bl[3955], bl[3956], bl[3957], bl[3958], bl[3959], bl[3960], bl[3961], bl[3962], bl[3963], bl[3964], bl[3965], bl[3966], bl[3967], bl[3968], bl[3969], bl[3970], bl[3971], bl[3972], bl[3973], bl[3974], bl[3975], bl[3976], bl[3977], bl[3978], bl[3979], bl[3980], bl[3981], bl[3982], bl[3983], bl[3984], bl[3985], bl[3986], bl[3987], bl[3988], bl[3989], bl[3990], bl[3991], bl[3992], bl[3993], bl[3994], bl[3995]}),
        .wl({wl[16], wl[17], wl[18], wl[19], wl[20], wl[21], wl[22], wl[23], wl[3996], wl[3997], wl[3998], wl[3999], wl[4000], wl[4001], wl[4002], wl[4003], wl[4004], wl[4005], wl[4006], wl[4007], wl[4008], wl[4009], wl[4010], wl[4011], wl[4012], wl[4013], wl[4014], wl[4015], wl[4016], wl[4017], wl[4018], wl[4019], wl[4020], wl[4021], wl[4022], wl[4023], wl[4024], wl[4025], wl[4026], wl[4027], wl[4028], wl[4029], wl[4030], wl[4031], wl[4032], wl[4033], wl[4034], wl[4035], wl[4036], wl[4037], wl[4038], wl[4039], wl[4040], wl[4041], wl[4042], wl[4043], wl[4044], wl[4045], wl[4046], wl[4047], wl[4048], wl[4049], wl[4050], wl[4051], wl[4052], wl[4053], wl[4054], wl[4055], wl[4056], wl[4057], wl[4058], wl[4059], wl[4060], wl[4061], wl[4062], wl[4063], wl[4064], wl[4065], wl[4066], wl[4067], wl[3918], wl[3919], wl[3920], wl[3921], wl[3922], wl[3923], wl[3924], wl[3925], wl[3926], wl[3927], wl[3928], wl[3929], wl[3930], wl[3931], wl[3932], wl[3933], wl[3934], wl[3935], wl[3936], wl[3937], wl[3938], wl[3939], wl[3940], wl[3941], wl[3942], wl[3943], wl[3944], wl[3945], wl[3946], wl[3947], wl[3948], wl[3949], wl[3950], wl[3951], wl[3952], wl[3953], wl[3954], wl[3955], wl[3956], wl[3957], wl[3958], wl[3959], wl[3960], wl[3961], wl[3962], wl[3963], wl[3964], wl[3965], wl[3966], wl[3967], wl[3968], wl[3969], wl[3970], wl[3971], wl[3972], wl[3973], wl[3974], wl[3975], wl[3976], wl[3977], wl[3978], wl[3979], wl[3980], wl[3981], wl[3982], wl[3983], wl[3984], wl[3985], wl[3986], wl[3987], wl[3988], wl[3989], wl[3990], wl[3991], wl[3992], wl[3993], wl[3994], wl[3995]})
    );
endmodule

