//Generated from netlist by SpyDrNet
//netlist name: SDN_VERILOG_NETLIST_logical_tile_io_mode_physical__iopad
module fpga_top
(
    reset,
    clk,
    gfpga_pad_GPIO_PAD
);

    input reset;
    input clk;
    inout [0:127]gfpga_pad_GPIO_PAD;

    wire reset;
    wire clk;
    wire [0:127]gfpga_pad_GPIO_PAD;
    wire [0:19]cbx_1__0__0_chanx_left_out;
    wire [0:19]cbx_1__0__0_chanx_right_out;
    wire [0:19]cbx_1__0__1_chanx_left_out;
    wire [0:19]cbx_1__0__1_chanx_right_out;
    wire [0:19]cbx_1__0__2_chanx_left_out;
    wire [0:19]cbx_1__0__2_chanx_right_out;
    wire [0:19]cbx_1__0__3_chanx_left_out;
    wire [0:19]cbx_1__0__3_chanx_right_out;
    wire [0:19]cbx_1__1__0_chanx_left_out;
    wire [0:19]cbx_1__1__0_chanx_right_out;
    wire [0:19]cbx_1__1__10_chanx_left_out;
    wire [0:19]cbx_1__1__10_chanx_right_out;
    wire [0:19]cbx_1__1__11_chanx_left_out;
    wire [0:19]cbx_1__1__11_chanx_right_out;
    wire [0:19]cbx_1__1__1_chanx_left_out;
    wire [0:19]cbx_1__1__1_chanx_right_out;
    wire [0:19]cbx_1__1__2_chanx_left_out;
    wire [0:19]cbx_1__1__2_chanx_right_out;
    wire [0:19]cbx_1__1__3_chanx_left_out;
    wire [0:19]cbx_1__1__3_chanx_right_out;
    wire [0:19]cbx_1__1__4_chanx_left_out;
    wire [0:19]cbx_1__1__4_chanx_right_out;
    wire [0:19]cbx_1__1__5_chanx_left_out;
    wire [0:19]cbx_1__1__5_chanx_right_out;
    wire [0:19]cbx_1__1__6_chanx_left_out;
    wire [0:19]cbx_1__1__6_chanx_right_out;
    wire [0:19]cbx_1__1__7_chanx_left_out;
    wire [0:19]cbx_1__1__7_chanx_right_out;
    wire [0:19]cbx_1__1__8_chanx_left_out;
    wire [0:19]cbx_1__1__8_chanx_right_out;
    wire [0:19]cbx_1__1__9_chanx_left_out;
    wire [0:19]cbx_1__1__9_chanx_right_out;
    wire [0:19]cbx_1__4__0_chanx_left_out;
    wire [0:19]cbx_1__4__0_chanx_right_out;
    wire [0:19]cbx_1__4__1_chanx_left_out;
    wire [0:19]cbx_1__4__1_chanx_right_out;
    wire [0:19]cbx_1__4__2_chanx_left_out;
    wire [0:19]cbx_1__4__2_chanx_right_out;
    wire [0:19]cbx_1__4__3_chanx_left_out;
    wire [0:19]cbx_1__4__3_chanx_right_out;
    wire [0:19]cby_0__1__0_chany_bottom_out;
    wire [0:19]cby_0__1__0_chany_top_out;
    wire [0:19]cby_0__1__1_chany_bottom_out;
    wire [0:19]cby_0__1__1_chany_top_out;
    wire [0:19]cby_0__1__2_chany_bottom_out;
    wire [0:19]cby_0__1__2_chany_top_out;
    wire [0:19]cby_0__1__3_chany_bottom_out;
    wire [0:19]cby_0__1__3_chany_top_out;
    wire [0:19]cby_1__1__0_chany_bottom_out;
    wire [0:19]cby_1__1__0_chany_top_out;
    wire [0:19]cby_1__1__10_chany_bottom_out;
    wire [0:19]cby_1__1__10_chany_top_out;
    wire [0:19]cby_1__1__11_chany_bottom_out;
    wire [0:19]cby_1__1__11_chany_top_out;
    wire [0:19]cby_1__1__1_chany_bottom_out;
    wire [0:19]cby_1__1__1_chany_top_out;
    wire [0:19]cby_1__1__2_chany_bottom_out;
    wire [0:19]cby_1__1__2_chany_top_out;
    wire [0:19]cby_1__1__3_chany_bottom_out;
    wire [0:19]cby_1__1__3_chany_top_out;
    wire [0:19]cby_1__1__4_chany_bottom_out;
    wire [0:19]cby_1__1__4_chany_top_out;
    wire [0:19]cby_1__1__5_chany_bottom_out;
    wire [0:19]cby_1__1__5_chany_top_out;
    wire [0:19]cby_1__1__6_chany_bottom_out;
    wire [0:19]cby_1__1__6_chany_top_out;
    wire [0:19]cby_1__1__7_chany_bottom_out;
    wire [0:19]cby_1__1__7_chany_top_out;
    wire [0:19]cby_1__1__8_chany_bottom_out;
    wire [0:19]cby_1__1__8_chany_top_out;
    wire [0:19]cby_1__1__9_chany_bottom_out;
    wire [0:19]cby_1__1__9_chany_top_out;
    wire [0:19]cby_4__1__0_chany_bottom_out;
    wire [0:19]cby_4__1__0_chany_top_out;
    wire [0:19]cby_4__1__1_chany_bottom_out;
    wire [0:19]cby_4__1__1_chany_top_out;
    wire [0:19]cby_4__1__2_chany_bottom_out;
    wire [0:19]cby_4__1__2_chany_top_out;
    wire [0:19]cby_4__1__3_chany_bottom_out;
    wire [0:19]cby_4__1__3_chany_top_out;
    wire [0:19]sb_0__0__0_chanx_right_out;
    wire [0:19]sb_0__0__0_chany_top_out;
    wire [0:19]sb_0__1__0_chanx_right_out;
    wire [0:19]sb_0__1__0_chany_bottom_out;
    wire [0:19]sb_0__1__0_chany_top_out;
    wire [0:19]sb_0__1__1_chanx_right_out;
    wire [0:19]sb_0__1__1_chany_bottom_out;
    wire [0:19]sb_0__1__1_chany_top_out;
    wire [0:19]sb_0__1__2_chanx_right_out;
    wire [0:19]sb_0__1__2_chany_bottom_out;
    wire [0:19]sb_0__1__2_chany_top_out;
    wire [0:19]sb_0__4__0_chanx_right_out;
    wire [0:19]sb_0__4__0_chany_bottom_out;
    wire [0:19]sb_1__0__0_chanx_left_out;
    wire [0:19]sb_1__0__0_chanx_right_out;
    wire [0:19]sb_1__0__0_chany_top_out;
    wire [0:19]sb_1__0__1_chanx_left_out;
    wire [0:19]sb_1__0__1_chanx_right_out;
    wire [0:19]sb_1__0__1_chany_top_out;
    wire [0:19]sb_1__0__2_chanx_left_out;
    wire [0:19]sb_1__0__2_chanx_right_out;
    wire [0:19]sb_1__0__2_chany_top_out;
    wire [0:19]sb_1__1__0_chanx_left_out;
    wire [0:19]sb_1__1__0_chanx_right_out;
    wire [0:19]sb_1__1__0_chany_bottom_out;
    wire [0:19]sb_1__1__0_chany_top_out;
    wire [0:19]sb_1__1__1_chanx_left_out;
    wire [0:19]sb_1__1__1_chanx_right_out;
    wire [0:19]sb_1__1__1_chany_bottom_out;
    wire [0:19]sb_1__1__1_chany_top_out;
    wire [0:19]sb_1__1__2_chanx_left_out;
    wire [0:19]sb_1__1__2_chanx_right_out;
    wire [0:19]sb_1__1__2_chany_bottom_out;
    wire [0:19]sb_1__1__2_chany_top_out;
    wire [0:19]sb_1__1__3_chanx_left_out;
    wire [0:19]sb_1__1__3_chanx_right_out;
    wire [0:19]sb_1__1__3_chany_bottom_out;
    wire [0:19]sb_1__1__3_chany_top_out;
    wire [0:19]sb_1__1__4_chanx_left_out;
    wire [0:19]sb_1__1__4_chanx_right_out;
    wire [0:19]sb_1__1__4_chany_bottom_out;
    wire [0:19]sb_1__1__4_chany_top_out;
    wire [0:19]sb_1__1__5_chanx_left_out;
    wire [0:19]sb_1__1__5_chanx_right_out;
    wire [0:19]sb_1__1__5_chany_bottom_out;
    wire [0:19]sb_1__1__5_chany_top_out;
    wire [0:19]sb_1__1__6_chanx_left_out;
    wire [0:19]sb_1__1__6_chanx_right_out;
    wire [0:19]sb_1__1__6_chany_bottom_out;
    wire [0:19]sb_1__1__6_chany_top_out;
    wire [0:19]sb_1__1__7_chanx_left_out;
    wire [0:19]sb_1__1__7_chanx_right_out;
    wire [0:19]sb_1__1__7_chany_bottom_out;
    wire [0:19]sb_1__1__7_chany_top_out;
    wire [0:19]sb_1__1__8_chanx_left_out;
    wire [0:19]sb_1__1__8_chanx_right_out;
    wire [0:19]sb_1__1__8_chany_bottom_out;
    wire [0:19]sb_1__1__8_chany_top_out;
    wire [0:19]sb_1__4__0_chanx_left_out;
    wire [0:19]sb_1__4__0_chanx_right_out;
    wire [0:19]sb_1__4__0_chany_bottom_out;
    wire [0:19]sb_1__4__1_chanx_left_out;
    wire [0:19]sb_1__4__1_chanx_right_out;
    wire [0:19]sb_1__4__1_chany_bottom_out;
    wire [0:19]sb_1__4__2_chanx_left_out;
    wire [0:19]sb_1__4__2_chanx_right_out;
    wire [0:19]sb_1__4__2_chany_bottom_out;
    wire [0:19]sb_4__0__0_chanx_left_out;
    wire [0:19]sb_4__0__0_chany_top_out;
    wire [0:19]sb_4__1__0_chanx_left_out;
    wire [0:19]sb_4__1__0_chany_bottom_out;
    wire [0:19]sb_4__1__0_chany_top_out;
    wire [0:19]sb_4__1__1_chanx_left_out;
    wire [0:19]sb_4__1__1_chany_bottom_out;
    wire [0:19]sb_4__1__1_chany_top_out;
    wire [0:19]sb_4__1__2_chanx_left_out;
    wire [0:19]sb_4__1__2_chany_bottom_out;
    wire [0:19]sb_4__1__2_chany_top_out;
    wire [0:19]sb_4__4__0_chanx_left_out;
    wire [0:19]sb_4__4__0_chany_bottom_out;
    wire [0:9]grid_clb_1__1__grid_left_in;
    wire [0:9]grid_clb_1__1__grid_top_in;
    wire [0:9]grid_clb_1__1__grid_right_in;
    wire [0:9]grid_clb_1__1__grid_bottom_in;
    wire [0:9]grid_clb_1__2__grid_left_in;
    wire [0:9]grid_clb_1__2__grid_top_in;
    wire [0:9]grid_clb_1__2__grid_right_in;
    wire [0:9]grid_clb_1__2__grid_bottom_in;
    wire [0:9]grid_clb_1__3__grid_left_in;
    wire [0:9]grid_clb_1__3__grid_top_in;
    wire [0:9]grid_clb_1__3__grid_right_in;
    wire [0:9]grid_clb_1__3__grid_bottom_in;
    wire [0:9]grid_clb_1__4__grid_left_in;
    wire [0:9]grid_clb_1__4__grid_top_in;
    wire [0:9]grid_clb_1__4__grid_right_in;
    wire [0:9]grid_clb_1__4__grid_bottom_in;
    wire [0:9]grid_clb_2__1__grid_left_in;
    wire [0:9]grid_clb_2__1__grid_top_in;
    wire [0:9]grid_clb_2__1__grid_right_in;
    wire [0:9]grid_clb_2__1__grid_bottom_in;
    wire [0:9]grid_clb_2__2__grid_left_in;
    wire [0:9]grid_clb_2__2__grid_top_in;
    wire [0:9]grid_clb_2__2__grid_right_in;
    wire [0:9]grid_clb_2__2__grid_bottom_in;
    wire [0:9]grid_clb_2__3__grid_left_in;
    wire [0:9]grid_clb_2__3__grid_top_in;
    wire [0:9]grid_clb_2__3__grid_right_in;
    wire [0:9]grid_clb_2__3__grid_bottom_in;
    wire [0:9]grid_clb_2__4__grid_left_in;
    wire [0:9]grid_clb_2__4__grid_top_in;
    wire [0:9]grid_clb_2__4__grid_right_in;
    wire [0:9]grid_clb_2__4__grid_bottom_in;
    wire [0:9]grid_clb_3__1__grid_left_in;
    wire [0:9]grid_clb_3__1__grid_top_in;
    wire [0:9]grid_clb_3__1__grid_right_in;
    wire [0:9]grid_clb_3__1__grid_bottom_in;
    wire [0:9]grid_clb_3__2__grid_left_in;
    wire [0:9]grid_clb_3__2__grid_top_in;
    wire [0:9]grid_clb_3__2__grid_right_in;
    wire [0:9]grid_clb_3__2__grid_bottom_in;
    wire [0:9]grid_clb_3__3__grid_left_in;
    wire [0:9]grid_clb_3__3__grid_top_in;
    wire [0:9]grid_clb_3__3__grid_right_in;
    wire [0:9]grid_clb_3__3__grid_bottom_in;
    wire [0:9]grid_clb_3__4__grid_left_in;
    wire [0:9]grid_clb_3__4__grid_top_in;
    wire [0:9]grid_clb_3__4__grid_right_in;
    wire [0:9]grid_clb_3__4__grid_bottom_in;
    wire [0:9]grid_clb_4__1__grid_left_in;
    wire [0:9]grid_clb_4__1__grid_top_in;
    wire [0:9]grid_clb_4__1__grid_right_in;
    wire [0:9]grid_clb_4__1__grid_bottom_in;
    wire [0:9]grid_clb_4__2__grid_left_in;
    wire [0:9]grid_clb_4__2__grid_top_in;
    wire [0:9]grid_clb_4__2__grid_right_in;
    wire [0:9]grid_clb_4__2__grid_bottom_in;
    wire [0:9]grid_clb_4__3__grid_left_in;
    wire [0:9]grid_clb_4__3__grid_top_in;
    wire [0:9]grid_clb_4__3__grid_right_in;
    wire [0:9]grid_clb_4__3__grid_bottom_in;
    wire [0:9]grid_clb_4__4__grid_left_in;
    wire [0:9]grid_clb_4__4__grid_top_in;
    wire [0:9]grid_clb_4__4__grid_right_in;
    wire [0:9]grid_clb_4__4__grid_bottom_in;
    wire [0:7]grid_io_top_1__5__io_bottom_in;
    wire [0:7]grid_io_top_1__5__io_bottom_out;
    wire [0:7]grid_io_top_2__5__io_bottom_in;
    wire [0:7]grid_io_top_2__5__io_bottom_out;
    wire [0:7]grid_io_top_3__5__io_bottom_in;
    wire [0:7]grid_io_top_3__5__io_bottom_out;
    wire [0:7]grid_io_top_4__5__io_bottom_in;
    wire [0:7]grid_io_top_4__5__io_bottom_out;
    wire [0:7]grid_io_right_5__4__io_left_in;
    wire [0:7]grid_io_right_5__4__io_left_out;
    wire [0:7]grid_io_right_5__3__io_left_in;
    wire [0:7]grid_io_right_5__3__io_left_out;
    wire [0:7]grid_io_right_5__2__io_left_in;
    wire [0:7]grid_io_right_5__2__io_left_out;
    wire [0:7]grid_io_right_5__1__io_left_in;
    wire [0:7]grid_io_right_5__1__io_left_out;
    wire [0:7]grid_io_bottom_4__0__io_top_in;
    wire [0:7]grid_io_bottom_4__0__io_top_out;
    wire [0:7]grid_io_bottom_3__0__io_top_in;
    wire [0:7]grid_io_bottom_3__0__io_top_out;
    wire [0:7]grid_io_bottom_2__0__io_top_in;
    wire [0:7]grid_io_bottom_2__0__io_top_out;
    wire [0:7]grid_io_bottom_1__0__io_top_in;
    wire [0:7]grid_io_bottom_1__0__io_top_out;
    wire [0:7]grid_io_left_0__1__io_right_in;
    wire [0:7]grid_io_left_0__1__io_right_out;
    wire [0:7]grid_io_left_0__2__io_right_in;
    wire [0:7]grid_io_left_0__2__io_right_out;
    wire [0:7]grid_io_left_0__3__io_right_in;
    wire [0:7]grid_io_left_0__3__io_right_out;
    wire [0:7]grid_io_left_0__4__io_right_in;
    wire [0:7]grid_io_left_0__4__io_right_out;
    wire [0:1]sb_0__0__grid_top_r_in;
    wire [0:1]sb_0__0__grid_right_t_in;
    wire [0:1]sb_0__1__grid_top_r_in;
    wire [0:1]sb_0__1__grid_right_t_in;
    wire [0:2]sb_0__1__grid_right_b_in;
    wire [0:1]sb_0__2__grid_top_r_in;
    wire [0:1]sb_0__2__grid_right_t_in;
    wire [0:2]sb_0__2__grid_right_b_in;
    wire [0:1]sb_0__3__grid_top_r_in;
    wire [0:1]sb_0__3__grid_right_t_in;
    wire [0:2]sb_0__3__grid_right_b_in;
    wire [0:2]sb_0__4__grid_right_b_in;
    wire [0:1]sb_1__0__grid_top_r_in;
    wire [0:2]sb_1__0__grid_top_l_in;
    wire [0:1]sb_1__0__grid_right_t_in;
    wire [0:1]sb_2__0__grid_top_r_in;
    wire [0:2]sb_2__0__grid_top_l_in;
    wire [0:1]sb_2__0__grid_right_t_in;
    wire [0:1]sb_3__0__grid_top_r_in;
    wire [0:2]sb_3__0__grid_top_l_in;
    wire [0:1]sb_3__0__grid_right_t_in;
    wire [0:1]sb_1__1__grid_top_r_in;
    wire [0:2]sb_1__1__grid_top_l_in;
    wire [0:1]sb_1__1__grid_right_t_in;
    wire [0:2]sb_1__1__grid_right_b_in;
    wire [0:1]sb_1__2__grid_top_r_in;
    wire [0:2]sb_1__2__grid_top_l_in;
    wire [0:1]sb_1__2__grid_right_t_in;
    wire [0:2]sb_1__2__grid_right_b_in;
    wire [0:1]sb_1__3__grid_top_r_in;
    wire [0:2]sb_1__3__grid_top_l_in;
    wire [0:1]sb_1__3__grid_right_t_in;
    wire [0:2]sb_1__3__grid_right_b_in;
    wire [0:1]sb_2__1__grid_top_r_in;
    wire [0:2]sb_2__1__grid_top_l_in;
    wire [0:1]sb_2__1__grid_right_t_in;
    wire [0:2]sb_2__1__grid_right_b_in;
    wire [0:1]sb_2__2__grid_top_r_in;
    wire [0:2]sb_2__2__grid_top_l_in;
    wire [0:1]sb_2__2__grid_right_t_in;
    wire [0:2]sb_2__2__grid_right_b_in;
    wire [0:1]sb_2__3__grid_top_r_in;
    wire [0:2]sb_2__3__grid_top_l_in;
    wire [0:1]sb_2__3__grid_right_t_in;
    wire [0:2]sb_2__3__grid_right_b_in;
    wire [0:1]sb_3__1__grid_top_r_in;
    wire [0:2]sb_3__1__grid_top_l_in;
    wire [0:1]sb_3__1__grid_right_t_in;
    wire [0:2]sb_3__1__grid_right_b_in;
    wire [0:1]sb_3__2__grid_top_r_in;
    wire [0:2]sb_3__2__grid_top_l_in;
    wire [0:1]sb_3__2__grid_right_t_in;
    wire [0:2]sb_3__2__grid_right_b_in;
    wire [0:1]sb_3__3__grid_top_r_in;
    wire [0:2]sb_3__3__grid_top_l_in;
    wire [0:1]sb_3__3__grid_right_t_in;
    wire [0:2]sb_3__3__grid_right_b_in;
    wire [0:2]sb_1__4__grid_right_b_in;
    wire [0:2]sb_2__4__grid_right_b_in;
    wire [0:2]sb_3__4__grid_right_b_in;
    wire [0:2]sb_4__0__grid_top_l_in;
    wire [0:2]sb_4__1__grid_top_l_in;
    wire [0:2]sb_4__2__grid_top_l_in;
    wire [0:2]sb_4__3__grid_top_l_in;

    tile tile_2__2_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_0__1__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_0__1__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_0__1__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_1__0__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_1__0__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_1__0__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_0__0__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_0__0__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_0__0__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_0__0__grid_top_r_in[1]),
        .grid_left_in(grid_clb_1__1__grid_left_in),
        .grid_bottom_in(grid_clb_1__1__grid_bottom_in),
        .chanx_left_in(sb_0__1__0_chanx_right_out),
        .chanx_left_out(cbx_1__1__0_chanx_left_out),
        .grid_top_out(grid_clb_1__2__grid_bottom_in),
        .chany_bottom_in(sb_1__0__0_chany_top_out),
        .chany_bottom_out(cby_1__1__0_chany_bottom_out),
        .grid_right_out(grid_clb_2__1__grid_left_in),
        .chany_top_in_0(cby_1__1__1_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__3_chanx_left_out),
        .chany_top_out_0(sb_1__1__0_chany_top_out),
        .chanx_right_out_0(sb_1__1__0_chanx_right_out),
        .grid_top_r_in(sb_1__1__grid_top_r_in),
        .grid_top_l_in(sb_1__1__grid_top_l_in),
        .grid_right_t_in(sb_1__1__grid_right_t_in),
        .grid_right_b_in(sb_1__1__grid_right_b_in),
        .grid_bottom_r_in(sb_1__0__grid_top_r_in),
        .grid_bottom_l_in(sb_1__0__grid_top_l_in),
        .grid_left_t_in(sb_0__1__grid_right_t_in),
        .grid_left_b_in(sb_0__1__grid_right_b_in),
        .bl({bl[1648], bl[1649], bl[1650], bl[1651], bl[1652], bl[1653], bl[1654], bl[1655], bl[1656], bl[1657], bl[1658], bl[1659], bl[1660], bl[1661], bl[1662], bl[1663], bl[1664], bl[1665], bl[1666], bl[1667], bl[1668], bl[1669], bl[1670], bl[1671], bl[1672], bl[1673], bl[1674], bl[1675], bl[1676], bl[1677], bl[1678], bl[1679], bl[1680], bl[1681], bl[1682], bl[1683], bl[1684], bl[1685], bl[1686], bl[1687], bl[1688], bl[1689], bl[1690], bl[1691], bl[1692], bl[1693], bl[1694], bl[1695], bl[1696], bl[1697], bl[1698], bl[1699], bl[1700], bl[1701], bl[1702], bl[1703], bl[1704], bl[1705], bl[1706], bl[1707], bl[1708], bl[1709], bl[1710], bl[1711], bl[1712], bl[1713], bl[1714], bl[1715], bl[1716], bl[1717], bl[1718], bl[1719], bl[1720], bl[1721], bl[1722], bl[1723], bl[1724], bl[1725], bl[1726], bl[1727], bl[1728], bl[1729], bl[1730], bl[1731], bl[1732], bl[1733], bl[1734], bl[1735], bl[1736], bl[1737], bl[1738], bl[1739], bl[1740], bl[1741], bl[1742], bl[1743], bl[1744], bl[1745], bl[1746], bl[1747], bl[1748], bl[1749], bl[1750], bl[1751], bl[1752], bl[1753], bl[1754], bl[1755], bl[1756], bl[1757], bl[1758], bl[1759], bl[1760], bl[1761], bl[1762], bl[1763], bl[1764], bl[1765], bl[1766], bl[1767], bl[1768], bl[1769], bl[1770], bl[1771], bl[1772], bl[1773], bl[1774], bl[1775], bl[1776], bl[1777], bl[1778], bl[1779], bl[1780], bl[1781], bl[1782], bl[1783], bl[1784], bl[1785], bl[1786], bl[1787], bl[1788], bl[1789], bl[1790], bl[1791], bl[1792], bl[1793], bl[1794], bl[1795], bl[1796], bl[1797], bl[1798], bl[1799], bl[1800], bl[1801], bl[1802], bl[1803], bl[1804], bl[1805], bl[1806], bl[1807], bl[1808], bl[1809], bl[1810], bl[1811], bl[1812], bl[1813], bl[1814], bl[1815], bl[1816], bl[1817], bl[1818], bl[1819], bl[1820], bl[1821], bl[1822], bl[1823], bl[1824], bl[1825], bl[1826], bl[1827], bl[1828], bl[1829], bl[1830], bl[1831], bl[1832], bl[1833], bl[1834], bl[1835], bl[1836], bl[1837], bl[1838], bl[1839], bl[1840], bl[1841], bl[1842], bl[1843], bl[1844], bl[1845], bl[1846], bl[1847], bl[1848], bl[1849], bl[1850], bl[1851], bl[1852], bl[1853], bl[1854], bl[1855], bl[1856], bl[1857], bl[1858], bl[1859], bl[1860], bl[1861], bl[1862], bl[1863], bl[1864], bl[1865], bl[1866], bl[1867], bl[1868], bl[1869], bl[1870], bl[1871], bl[1872], bl[1873], bl[1874], bl[1875], bl[1876], bl[1877], bl[1878], bl[1879], bl[1880], bl[1881], bl[1882], bl[1883], bl[1884], bl[1885], bl[1886], bl[1887], bl[1888], bl[1889], bl[1890], bl[1891], bl[1892], bl[1893], bl[1894], bl[1895], bl[1896], bl[1897], bl[1898], bl[1899], bl[1900], bl[1901], bl[1902], bl[1903], bl[1904], bl[1905], bl[1906], bl[1907], bl[1908], bl[1909], bl[1910], bl[1911], bl[1912], bl[1913], bl[1914], bl[1915], bl[1916], bl[1917], bl[1918], bl[1919], bl[1920], bl[1921], bl[1922], bl[1923], bl[1924], bl[1925], bl[1926], bl[1927], bl[1928], bl[1929], bl[1930], bl[1931], bl[1932], bl[1933], bl[1934], bl[1935], bl[1936], bl[1937], bl[1938], bl[1939], bl[1940], bl[1941], bl[1942], bl[1943], bl[1944], bl[1945], bl[1946], bl[1947], bl[1948], bl[1949], bl[1950], bl[1951], bl[1952], bl[1953], bl[1954], bl[1955], bl[1956], bl[1957], bl[1958], bl[1959], bl[1960], bl[1961], bl[1962], bl[1963], bl[1964], bl[1965], bl[1966], bl[1967], bl[1968], bl[1969], bl[1970], bl[1971], bl[1972], bl[1973], bl[1974], bl[1975], bl[1976], bl[1977], bl[1978], bl[1979], bl[1980], bl[1981], bl[1982], bl[1983], bl[1984], bl[1985], bl[1986], bl[1987], bl[1988], bl[1989], bl[1990], bl[1991], bl[1992], bl[1993], bl[1994], bl[1995], bl[1996], bl[1997], bl[1998], bl[1999], bl[2000], bl[2001], bl[2002], bl[2003], bl[2004], bl[2005], bl[2006], bl[2007], bl[2008], bl[2009], bl[2010], bl[2011], bl[2012], bl[2013], bl[2014], bl[2015], bl[2016], bl[2017], bl[2018], bl[2019], bl[2020], bl[2021], bl[2022], bl[2023], bl[2024], bl[2025], bl[2026], bl[2027], bl[2028], bl[2029], bl[2030], bl[2031], bl[2032], bl[2033], bl[2034], bl[2035], bl[2036], bl[2037], bl[2038], bl[2039], bl[2040], bl[2041], bl[2042], bl[2043], bl[2044], bl[2045], bl[2046], bl[2047], bl[2048], bl[2049], bl[2050], bl[2051], bl[2052], bl[2053], bl[2054], bl[2055], bl[2056], bl[2057], bl[2058], bl[2059], bl[2060], bl[2061], bl[2062], bl[2063], bl[2064], bl[2065], bl[2066], bl[2067], bl[2068], bl[2069], bl[2070], bl[2071], bl[2072], bl[2073], bl[2074], bl[2075], bl[2076], bl[2077], bl[2078], bl[2079], bl[2080], bl[2081], bl[2082], bl[2083], bl[2084], bl[2085], bl[2086], bl[2087], bl[2088], bl[2089], bl[2090], bl[2091], bl[2092], bl[2093], bl[2094], bl[2095], bl[2096], bl[2097], bl[2098], bl[2099], bl[2100], bl[2101], bl[2102], bl[2103], bl[2104], bl[2105], bl[2106], bl[2107], bl[2108], bl[2109], bl[2110], bl[2111], bl[2112], bl[2113], bl[2114], bl[2115], bl[2116], bl[2117], bl[2118], bl[2119], bl[2120], bl[2121], bl[2122], bl[2123], bl[2124], bl[2125], bl[2126], bl[2127], bl[2128], bl[2129], bl[2130], bl[2131], bl[2132], bl[2133], bl[2134], bl[2135], bl[2136], bl[2137], bl[2138], bl[2139], bl[2140], bl[2141], bl[2142], bl[2143], bl[2144], bl[2145], bl[2146], bl[2147], bl[2148], bl[2149], bl[2150], bl[2151], bl[2152], bl[2153], bl[2154], bl[2155], bl[2156], bl[2157], bl[2158], bl[2159], bl[2160], bl[2161], bl[2162], bl[2163], bl[2164], bl[2165], bl[2166], bl[2167], bl[2168], bl[2169], bl[2170], bl[2171], bl[2172], bl[2173], bl[2174], bl[2175], bl[2176], bl[2177], bl[2178], bl[2179], bl[2180], bl[2181], bl[2182], bl[2183], bl[2184], bl[2185], bl[2186], bl[2187], bl[2188], bl[2189], bl[2190], bl[2191], bl[2192], bl[2193], bl[2194], bl[2195], bl[2196], bl[2197], bl[2198], bl[2199], bl[2200], bl[2201], bl[2202], bl[2203], bl[2204], bl[2205], bl[2206], bl[2207], bl[2208], bl[2209], bl[2210], bl[2211], bl[2212], bl[2213], bl[2214], bl[2215], bl[2216], bl[2217], bl[2218], bl[2219], bl[2220], bl[2221], bl[2222], bl[2223], bl[2224], bl[2225], bl[2226], bl[2227], bl[2228], bl[2229], bl[2230], bl[2231], bl[2232], bl[2233], bl[2234], bl[2235], bl[2236], bl[2237], bl[2238], bl[2239], bl[2240], bl[2241], bl[2242], bl[2243], bl[2244], bl[2245], bl[2246], bl[2247], bl[2248], bl[2249], bl[2250], bl[2251], bl[2252], bl[2253], bl[2254], bl[2255], bl[2256], bl[2257], bl[2258], bl[2259], bl[2260], bl[2261], bl[2262], bl[2263], bl[2264], bl[2265], bl[2266], bl[2267], bl[2268], bl[2269], bl[2270], bl[2271], bl[2272], bl[2273], bl[2274], bl[2275], bl[2276], bl[2277], bl[2278], bl[2279], bl[2280], bl[2281], bl[2282], bl[2283], bl[2284], bl[2285], bl[2286], bl[2287], bl[2288], bl[2289], bl[2290], bl[2291], bl[2292], bl[2293], bl[2294], bl[2295], bl[2296], bl[2297], bl[2298], bl[2299], bl[2300], bl[2301], bl[2302], bl[2303], bl[2304], bl[2305], bl[2306], bl[2307], bl[2308], bl[2309], bl[2310], bl[2311], bl[2312], bl[2313], bl[2314], bl[2315], bl[2316], bl[2317], bl[2318], bl[2319], bl[2320], bl[2321], bl[2322], bl[2323], bl[2324], bl[2325], bl[2326], bl[2327], bl[2328], bl[2329], bl[2330], bl[2331], bl[2332], bl[2333], bl[2334], bl[2335], bl[2336], bl[2337], bl[2338], bl[2339], bl[2340], bl[2341], bl[2342], bl[2343], bl[2344], bl[2345], bl[2346], bl[2347], bl[2348], bl[2349], bl[2350], bl[2351], bl[2352], bl[2353], bl[2354], bl[2355], bl[2356], bl[2357], bl[2358], bl[2359], bl[2360], bl[2361], bl[2362], bl[2363], bl[2364], bl[2365], bl[2366], bl[2367], bl[2368], bl[2369], bl[2370], bl[2371], bl[2372], bl[2373], bl[2374], bl[2375], bl[2376], bl[2377], bl[2378], bl[2379], bl[2380], bl[2381], bl[2382], bl[2383], bl[2384], bl[2385], bl[2386], bl[2387], bl[2388], bl[2389], bl[2390], bl[2391], bl[2392], bl[2393], bl[2394], bl[2395], bl[2396], bl[2397], bl[2398], bl[2399], bl[2400], bl[2401], bl[2402], bl[2403], bl[2404], bl[2405], bl[2406], bl[2407], bl[2408], bl[2409], bl[2410], bl[2411], bl[2412], bl[2413], bl[2414], bl[2415], bl[2416], bl[2417], bl[2418], bl[2419], bl[2420], bl[2421], bl[2422], bl[2423], bl[2424], bl[2425], bl[2426], bl[2427], bl[2428], bl[2429], bl[2430], bl[2431], bl[2432], bl[2433], bl[2434], bl[2435], bl[2436], bl[2437], bl[2438], bl[2439], bl[2440], bl[2441], bl[2442], bl[2443], bl[2444], bl[2445], bl[2446], bl[2447], bl[2448], bl[2449], bl[2450], bl[2451], bl[2452], bl[2453], bl[2454], bl[2455], bl[2456], bl[2457], bl[2458], bl[2459], bl[2460], bl[2461], bl[2462], bl[2463], bl[2464], bl[2465], bl[2466], bl[2467], bl[2468], bl[2469], bl[2470], bl[2471], bl[2472], bl[2473], bl[2474], bl[2475], bl[2476], bl[2477], bl[2478], bl[2479], bl[2480], bl[2481], bl[2482], bl[2483], bl[2484], bl[2485], bl[2486], bl[2487], bl[2488], bl[2489], bl[2490], bl[2491], bl[2492], bl[2493], bl[2494], bl[2495], bl[2496], bl[2497], bl[2498], bl[2499], bl[2500], bl[2501], bl[2502], bl[2503], bl[2504], bl[2505], bl[2506], bl[2507], bl[2508], bl[2509], bl[2510], bl[2511], bl[2512], bl[2513], bl[2514], bl[2515], bl[2516], bl[2517], bl[2518], bl[2519], bl[2520], bl[2521], bl[2522], bl[2523], bl[2524], bl[2525], bl[2526], bl[2527], bl[2528], bl[2529], bl[2530], bl[2531], bl[2532], bl[2533], bl[2534], bl[2535], bl[2536], bl[2537], bl[2538], bl[2539], bl[2540], bl[2541], bl[2542], bl[2543], bl[2544], bl[2545], bl[2546], bl[2547], bl[2548], bl[2549], bl[2550], bl[2551], bl[2552], bl[2553], bl[2554], bl[2555], bl[2556], bl[2557], bl[2558], bl[2559], bl[2560], bl[2561], bl[2562], bl[2563], bl[2564], bl[2565], bl[2566], bl[2567], bl[2568], bl[2569], bl[2570], bl[2571], bl[2572], bl[2573], bl[2574], bl[2575], bl[2576], bl[2577], bl[2578], bl[2579], bl[2580], bl[2581], bl[2582], bl[2583], bl[2584], bl[2585], bl[2586], bl[2587], bl[2588], bl[2589], bl[2590], bl[2591], bl[2592], bl[2593], bl[2594], bl[2595], bl[2596], bl[2597], bl[2598], bl[2599], bl[2600], bl[2601], bl[2602], bl[2603], bl[2604], bl[2605], bl[2606], bl[2607], bl[2608], bl[2609], bl[2610], bl[2611], bl[2612], bl[2613], bl[2614], bl[2615], bl[2616], bl[2617], bl[2618], bl[2619], bl[2620], bl[2621], bl[2622], bl[2623], bl[2624], bl[2625], bl[2626], bl[2627], bl[2628], bl[2629], bl[2630], bl[2631], bl[2632], bl[2633], bl[2634], bl[2635], bl[2636], bl[2637], bl[2638], bl[2639], bl[2640], bl[2641], bl[2642], bl[2643], bl[2644], bl[2645], bl[2646], bl[2647], bl[2648], bl[2649], bl[2650], bl[2651], bl[2652], bl[2653], bl[2654], bl[2655], bl[2656], bl[2657], bl[2658], bl[2659], bl[2660], bl[2661], bl[2662], bl[2663], bl[2664], bl[2665], bl[2666], bl[2667], bl[10264], bl[10265], bl[10266], bl[10267], bl[10268], bl[10269], bl[10270], bl[10271], bl[10272], bl[10273], bl[10274], bl[10275], bl[10276], bl[10277], bl[10278], bl[10279], bl[10280], bl[10281], bl[10282], bl[10283], bl[10284], bl[10285], bl[10286], bl[10287], bl[10288], bl[10289], bl[10290], bl[10291], bl[10292], bl[10293], bl[10294], bl[10295], bl[10296], bl[10297], bl[10298], bl[10299], bl[10300], bl[10301], bl[10302], bl[10303], bl[10304], bl[10305], bl[10306], bl[10307], bl[10308], bl[10309], bl[10310], bl[10311], bl[10312], bl[10313], bl[10314], bl[10315], bl[10316], bl[10317], bl[10318], bl[10319], bl[10320], bl[10321], bl[10322], bl[10323], bl[10324], bl[10325], bl[10326], bl[10327], bl[10328], bl[10329], bl[10330], bl[10331], bl[10332], bl[10333], bl[10334], bl[10335], bl[10336], bl[10337], bl[10338], bl[10339], bl[10340], bl[10341], bl[10342], bl[10343], bl[1568], bl[1569], bl[1570], bl[1571], bl[1572], bl[1573], bl[1574], bl[1575], bl[1576], bl[1577], bl[1578], bl[1579], bl[1580], bl[1581], bl[1582], bl[1583], bl[1584], bl[1585], bl[1586], bl[1587], bl[1588], bl[1589], bl[1590], bl[1591], bl[1592], bl[1593], bl[1594], bl[1595], bl[1596], bl[1597], bl[1598], bl[1599], bl[1600], bl[1601], bl[1602], bl[1603], bl[1604], bl[1605], bl[1606], bl[1607], bl[1608], bl[1609], bl[1610], bl[1611], bl[1612], bl[1613], bl[1614], bl[1615], bl[1616], bl[1617], bl[1618], bl[1619], bl[1620], bl[1621], bl[1622], bl[1623], bl[1624], bl[1625], bl[1626], bl[1627], bl[1628], bl[1629], bl[1630], bl[1631], bl[1632], bl[1633], bl[1634], bl[1635], bl[1636], bl[1637], bl[1638], bl[1639], bl[1640], bl[1641], bl[1642], bl[1643], bl[1644], bl[1645], bl[1646], bl[1647], bl[10184], bl[10185], bl[10186], bl[10187], bl[10188], bl[10189], bl[10190], bl[10191], bl[10192], bl[10193], bl[10194], bl[10195], bl[10196], bl[10197], bl[10198], bl[10199], bl[10200], bl[10201], bl[10202], bl[10203], bl[10204], bl[10205], bl[10206], bl[10207], bl[10208], bl[10209], bl[10210], bl[10211], bl[10212], bl[10213], bl[10214], bl[10215], bl[10216], bl[10217], bl[10218], bl[10219], bl[10220], bl[10221], bl[10222], bl[10223], bl[10224], bl[10225], bl[10226], bl[10227], bl[10228], bl[10229], bl[10230], bl[10231], bl[10232], bl[10233], bl[10234], bl[10235], bl[10236], bl[10237], bl[10238], bl[10239], bl[10240], bl[10241], bl[10242], bl[10243], bl[10244], bl[10245], bl[10246], bl[10247], bl[10248], bl[10249], bl[10250], bl[10251], bl[10252], bl[10253], bl[10254], bl[10255], bl[10256], bl[10257], bl[10258], bl[10259], bl[10260], bl[10261], bl[10262], bl[10263]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    tile tile_2__3_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_0__2__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_0__2__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_0__2__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_1__1__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_1__1__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_1__1__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_0__1__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_0__1__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_0__1__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_0__1__grid_top_r_in[1]),
        .grid_left_in(grid_clb_1__2__grid_left_in),
        .grid_bottom_in(grid_clb_1__2__grid_bottom_in),
        .chanx_left_in(sb_0__1__1_chanx_right_out),
        .chanx_left_out(cbx_1__1__1_chanx_left_out),
        .grid_top_out(grid_clb_1__3__grid_bottom_in),
        .chany_bottom_in(sb_1__1__0_chany_top_out),
        .chany_bottom_out(cby_1__1__1_chany_bottom_out),
        .grid_right_out(grid_clb_2__2__grid_left_in),
        .chany_top_in_0(cby_1__1__2_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__4_chanx_left_out),
        .chany_top_out_0(sb_1__1__1_chany_top_out),
        .chanx_right_out_0(sb_1__1__1_chanx_right_out),
        .grid_top_r_in(sb_1__2__grid_top_r_in),
        .grid_top_l_in(sb_1__2__grid_top_l_in),
        .grid_right_t_in(sb_1__2__grid_right_t_in),
        .grid_right_b_in(sb_1__2__grid_right_b_in),
        .grid_bottom_r_in(sb_1__1__grid_top_r_in),
        .grid_bottom_l_in(sb_1__1__grid_top_l_in),
        .grid_left_t_in(sb_0__2__grid_right_t_in),
        .grid_left_b_in(sb_0__2__grid_right_b_in),
        .bl({bl[10424], bl[10425], bl[10426], bl[10427], bl[10428], bl[10429], bl[10430], bl[10431], bl[10432], bl[10433], bl[10434], bl[10435], bl[10436], bl[10437], bl[10438], bl[10439], bl[10440], bl[10441], bl[10442], bl[10443], bl[10444], bl[10445], bl[10446], bl[10447], bl[10448], bl[10449], bl[10450], bl[10451], bl[10452], bl[10453], bl[10454], bl[10455], bl[10456], bl[10457], bl[10458], bl[10459], bl[10460], bl[10461], bl[10462], bl[10463], bl[10464], bl[10465], bl[10466], bl[10467], bl[10468], bl[10469], bl[10470], bl[10471], bl[10472], bl[10473], bl[10474], bl[10475], bl[10476], bl[10477], bl[10478], bl[10479], bl[10480], bl[10481], bl[10482], bl[10483], bl[10484], bl[10485], bl[10486], bl[10487], bl[10488], bl[10489], bl[10490], bl[10491], bl[10492], bl[10493], bl[10494], bl[10495], bl[10496], bl[10497], bl[10498], bl[10499], bl[10500], bl[10501], bl[10502], bl[10503], bl[10504], bl[10505], bl[10506], bl[10507], bl[10508], bl[10509], bl[10510], bl[10511], bl[10512], bl[10513], bl[10514], bl[10515], bl[10516], bl[10517], bl[10518], bl[10519], bl[10520], bl[10521], bl[10522], bl[10523], bl[10524], bl[10525], bl[10526], bl[10527], bl[10528], bl[10529], bl[10530], bl[10531], bl[10532], bl[10533], bl[10534], bl[10535], bl[10536], bl[10537], bl[10538], bl[10539], bl[10540], bl[10541], bl[10542], bl[10543], bl[10544], bl[10545], bl[10546], bl[10547], bl[10548], bl[10549], bl[10550], bl[10551], bl[10552], bl[10553], bl[10554], bl[10555], bl[10556], bl[10557], bl[10558], bl[10559], bl[10560], bl[10561], bl[10562], bl[10563], bl[10564], bl[10565], bl[10566], bl[10567], bl[10568], bl[10569], bl[10570], bl[10571], bl[10572], bl[10573], bl[10574], bl[10575], bl[10576], bl[10577], bl[10578], bl[10579], bl[10580], bl[10581], bl[10582], bl[10583], bl[10584], bl[10585], bl[10586], bl[10587], bl[10588], bl[10589], bl[10590], bl[10591], bl[10592], bl[10593], bl[10594], bl[10595], bl[10596], bl[10597], bl[10598], bl[10599], bl[10600], bl[10601], bl[10602], bl[10603], bl[10604], bl[10605], bl[10606], bl[10607], bl[10608], bl[10609], bl[10610], bl[10611], bl[10612], bl[10613], bl[10614], bl[10615], bl[10616], bl[10617], bl[10618], bl[10619], bl[10620], bl[10621], bl[10622], bl[10623], bl[10624], bl[10625], bl[10626], bl[10627], bl[10628], bl[10629], bl[10630], bl[10631], bl[10632], bl[10633], bl[10634], bl[10635], bl[10636], bl[10637], bl[10638], bl[10639], bl[10640], bl[10641], bl[10642], bl[10643], bl[10644], bl[10645], bl[10646], bl[10647], bl[10648], bl[10649], bl[10650], bl[10651], bl[10652], bl[10653], bl[10654], bl[10655], bl[10656], bl[10657], bl[10658], bl[10659], bl[10660], bl[10661], bl[10662], bl[10663], bl[10664], bl[10665], bl[10666], bl[10667], bl[10668], bl[10669], bl[10670], bl[10671], bl[10672], bl[10673], bl[10674], bl[10675], bl[10676], bl[10677], bl[10678], bl[10679], bl[10680], bl[10681], bl[10682], bl[10683], bl[10684], bl[10685], bl[10686], bl[10687], bl[10688], bl[10689], bl[10690], bl[10691], bl[10692], bl[10693], bl[10694], bl[10695], bl[10696], bl[10697], bl[10698], bl[10699], bl[10700], bl[10701], bl[10702], bl[10703], bl[10704], bl[10705], bl[10706], bl[10707], bl[10708], bl[10709], bl[10710], bl[10711], bl[10712], bl[10713], bl[10714], bl[10715], bl[10716], bl[10717], bl[10718], bl[10719], bl[10720], bl[10721], bl[10722], bl[10723], bl[10724], bl[10725], bl[10726], bl[10727], bl[10728], bl[10729], bl[10730], bl[10731], bl[10732], bl[10733], bl[10734], bl[10735], bl[10736], bl[10737], bl[10738], bl[10739], bl[10740], bl[10741], bl[10742], bl[10743], bl[10744], bl[10745], bl[10746], bl[10747], bl[10748], bl[10749], bl[10750], bl[10751], bl[10752], bl[10753], bl[10754], bl[10755], bl[10756], bl[10757], bl[10758], bl[10759], bl[10760], bl[10761], bl[10762], bl[10763], bl[10764], bl[10765], bl[10766], bl[10767], bl[10768], bl[10769], bl[10770], bl[10771], bl[10772], bl[10773], bl[10774], bl[10775], bl[10776], bl[10777], bl[10778], bl[10779], bl[10780], bl[10781], bl[10782], bl[10783], bl[10784], bl[10785], bl[10786], bl[10787], bl[10788], bl[10789], bl[10790], bl[10791], bl[10792], bl[10793], bl[10794], bl[10795], bl[10796], bl[10797], bl[10798], bl[10799], bl[10800], bl[10801], bl[10802], bl[10803], bl[10804], bl[10805], bl[10806], bl[10807], bl[10808], bl[10809], bl[10810], bl[10811], bl[10812], bl[10813], bl[10814], bl[10815], bl[10816], bl[10817], bl[10818], bl[10819], bl[10820], bl[10821], bl[10822], bl[10823], bl[10824], bl[10825], bl[10826], bl[10827], bl[10828], bl[10829], bl[10830], bl[10831], bl[10832], bl[10833], bl[10834], bl[10835], bl[10836], bl[10837], bl[10838], bl[10839], bl[10840], bl[10841], bl[10842], bl[10843], bl[10844], bl[10845], bl[10846], bl[10847], bl[10848], bl[10849], bl[10850], bl[10851], bl[10852], bl[10853], bl[10854], bl[10855], bl[10856], bl[10857], bl[10858], bl[10859], bl[10860], bl[10861], bl[10862], bl[10863], bl[10864], bl[10865], bl[10866], bl[10867], bl[10868], bl[10869], bl[10870], bl[10871], bl[10872], bl[10873], bl[10874], bl[10875], bl[10876], bl[10877], bl[10878], bl[10879], bl[10880], bl[10881], bl[10882], bl[10883], bl[10884], bl[10885], bl[10886], bl[10887], bl[10888], bl[10889], bl[10890], bl[10891], bl[10892], bl[10893], bl[10894], bl[10895], bl[10896], bl[10897], bl[10898], bl[10899], bl[10900], bl[10901], bl[10902], bl[10903], bl[10904], bl[10905], bl[10906], bl[10907], bl[10908], bl[10909], bl[10910], bl[10911], bl[10912], bl[10913], bl[10914], bl[10915], bl[10916], bl[10917], bl[10918], bl[10919], bl[10920], bl[10921], bl[10922], bl[10923], bl[10924], bl[10925], bl[10926], bl[10927], bl[10928], bl[10929], bl[10930], bl[10931], bl[10932], bl[10933], bl[10934], bl[10935], bl[10936], bl[10937], bl[10938], bl[10939], bl[10940], bl[10941], bl[10942], bl[10943], bl[10944], bl[10945], bl[10946], bl[10947], bl[10948], bl[10949], bl[10950], bl[10951], bl[10952], bl[10953], bl[10954], bl[10955], bl[10956], bl[10957], bl[10958], bl[10959], bl[10960], bl[10961], bl[10962], bl[10963], bl[10964], bl[10965], bl[10966], bl[10967], bl[10968], bl[10969], bl[10970], bl[10971], bl[10972], bl[10973], bl[10974], bl[10975], bl[10976], bl[10977], bl[10978], bl[10979], bl[10980], bl[10981], bl[10982], bl[10983], bl[10984], bl[10985], bl[10986], bl[10987], bl[10988], bl[10989], bl[10990], bl[10991], bl[10992], bl[10993], bl[10994], bl[10995], bl[10996], bl[10997], bl[10998], bl[10999], bl[11000], bl[11001], bl[11002], bl[11003], bl[11004], bl[11005], bl[11006], bl[11007], bl[11008], bl[11009], bl[11010], bl[11011], bl[11012], bl[11013], bl[11014], bl[11015], bl[11016], bl[11017], bl[11018], bl[11019], bl[11020], bl[11021], bl[11022], bl[11023], bl[11024], bl[11025], bl[11026], bl[11027], bl[11028], bl[11029], bl[11030], bl[11031], bl[11032], bl[11033], bl[11034], bl[11035], bl[11036], bl[11037], bl[11038], bl[11039], bl[11040], bl[11041], bl[11042], bl[11043], bl[11044], bl[11045], bl[11046], bl[11047], bl[11048], bl[11049], bl[11050], bl[11051], bl[11052], bl[11053], bl[11054], bl[11055], bl[11056], bl[11057], bl[11058], bl[11059], bl[11060], bl[11061], bl[11062], bl[11063], bl[11064], bl[11065], bl[11066], bl[11067], bl[11068], bl[11069], bl[11070], bl[11071], bl[11072], bl[11073], bl[11074], bl[11075], bl[11076], bl[11077], bl[11078], bl[11079], bl[11080], bl[11081], bl[11082], bl[11083], bl[11084], bl[11085], bl[11086], bl[11087], bl[11088], bl[11089], bl[11090], bl[11091], bl[11092], bl[11093], bl[11094], bl[11095], bl[11096], bl[11097], bl[11098], bl[11099], bl[11100], bl[11101], bl[11102], bl[11103], bl[11104], bl[11105], bl[11106], bl[11107], bl[11108], bl[11109], bl[11110], bl[11111], bl[11112], bl[11113], bl[11114], bl[11115], bl[11116], bl[11117], bl[11118], bl[11119], bl[11120], bl[11121], bl[11122], bl[11123], bl[11124], bl[11125], bl[11126], bl[11127], bl[11128], bl[11129], bl[11130], bl[11131], bl[11132], bl[11133], bl[11134], bl[11135], bl[11136], bl[11137], bl[11138], bl[11139], bl[11140], bl[11141], bl[11142], bl[11143], bl[11144], bl[11145], bl[11146], bl[11147], bl[11148], bl[11149], bl[11150], bl[11151], bl[11152], bl[11153], bl[11154], bl[11155], bl[11156], bl[11157], bl[11158], bl[11159], bl[11160], bl[11161], bl[11162], bl[11163], bl[11164], bl[11165], bl[11166], bl[11167], bl[11168], bl[11169], bl[11170], bl[11171], bl[11172], bl[11173], bl[11174], bl[11175], bl[11176], bl[11177], bl[11178], bl[11179], bl[11180], bl[11181], bl[11182], bl[11183], bl[11184], bl[11185], bl[11186], bl[11187], bl[11188], bl[11189], bl[11190], bl[11191], bl[11192], bl[11193], bl[11194], bl[11195], bl[11196], bl[11197], bl[11198], bl[11199], bl[11200], bl[11201], bl[11202], bl[11203], bl[11204], bl[11205], bl[11206], bl[11207], bl[11208], bl[11209], bl[11210], bl[11211], bl[11212], bl[11213], bl[11214], bl[11215], bl[11216], bl[11217], bl[11218], bl[11219], bl[11220], bl[11221], bl[11222], bl[11223], bl[11224], bl[11225], bl[11226], bl[11227], bl[11228], bl[11229], bl[11230], bl[11231], bl[11232], bl[11233], bl[11234], bl[11235], bl[11236], bl[11237], bl[11238], bl[11239], bl[11240], bl[11241], bl[11242], bl[11243], bl[11244], bl[11245], bl[11246], bl[11247], bl[11248], bl[11249], bl[11250], bl[11251], bl[11252], bl[11253], bl[11254], bl[11255], bl[11256], bl[11257], bl[11258], bl[11259], bl[11260], bl[11261], bl[11262], bl[11263], bl[11264], bl[11265], bl[11266], bl[11267], bl[11268], bl[11269], bl[11270], bl[11271], bl[11272], bl[11273], bl[11274], bl[11275], bl[11276], bl[11277], bl[11278], bl[11279], bl[11280], bl[11281], bl[11282], bl[11283], bl[11284], bl[11285], bl[11286], bl[11287], bl[11288], bl[11289], bl[11290], bl[11291], bl[11292], bl[11293], bl[11294], bl[11295], bl[11296], bl[11297], bl[11298], bl[11299], bl[11300], bl[11301], bl[11302], bl[11303], bl[11304], bl[11305], bl[11306], bl[11307], bl[11308], bl[11309], bl[11310], bl[11311], bl[11312], bl[11313], bl[11314], bl[11315], bl[11316], bl[11317], bl[11318], bl[11319], bl[11320], bl[11321], bl[11322], bl[11323], bl[11324], bl[11325], bl[11326], bl[11327], bl[11328], bl[11329], bl[11330], bl[11331], bl[11332], bl[11333], bl[11334], bl[11335], bl[11336], bl[11337], bl[11338], bl[11339], bl[11340], bl[11341], bl[11342], bl[11343], bl[11344], bl[11345], bl[11346], bl[11347], bl[11348], bl[11349], bl[11350], bl[11351], bl[11352], bl[11353], bl[11354], bl[11355], bl[11356], bl[11357], bl[11358], bl[11359], bl[11360], bl[11361], bl[11362], bl[11363], bl[11364], bl[11365], bl[11366], bl[11367], bl[11368], bl[11369], bl[11370], bl[11371], bl[11372], bl[11373], bl[11374], bl[11375], bl[11376], bl[11377], bl[11378], bl[11379], bl[11380], bl[11381], bl[11382], bl[11383], bl[11384], bl[11385], bl[11386], bl[11387], bl[11388], bl[11389], bl[11390], bl[11391], bl[11392], bl[11393], bl[11394], bl[11395], bl[11396], bl[11397], bl[11398], bl[11399], bl[11400], bl[11401], bl[11402], bl[11403], bl[11404], bl[11405], bl[11406], bl[11407], bl[11408], bl[11409], bl[11410], bl[11411], bl[11412], bl[11413], bl[11414], bl[11415], bl[11416], bl[11417], bl[11418], bl[11419], bl[11420], bl[11421], bl[11422], bl[11423], bl[11424], bl[11425], bl[11426], bl[11427], bl[11428], bl[11429], bl[11430], bl[11431], bl[11432], bl[11433], bl[11434], bl[11435], bl[11436], bl[11437], bl[11438], bl[11439], bl[11440], bl[11441], bl[11442], bl[11443], bl[11524], bl[11525], bl[11526], bl[11527], bl[11528], bl[11529], bl[11530], bl[11531], bl[11532], bl[11533], bl[11534], bl[11535], bl[11536], bl[11537], bl[11538], bl[11539], bl[11540], bl[11541], bl[11542], bl[11543], bl[11544], bl[11545], bl[11546], bl[11547], bl[11548], bl[11549], bl[11550], bl[11551], bl[11552], bl[11553], bl[11554], bl[11555], bl[11556], bl[11557], bl[11558], bl[11559], bl[11560], bl[11561], bl[11562], bl[11563], bl[11564], bl[11565], bl[11566], bl[11567], bl[11568], bl[11569], bl[11570], bl[11571], bl[11572], bl[11573], bl[11574], bl[11575], bl[11576], bl[11577], bl[11578], bl[11579], bl[11580], bl[11581], bl[11582], bl[11583], bl[11584], bl[11585], bl[11586], bl[11587], bl[11588], bl[11589], bl[11590], bl[11591], bl[11592], bl[11593], bl[11594], bl[11595], bl[11596], bl[11597], bl[11598], bl[11599], bl[11600], bl[11601], bl[11602], bl[11603], bl[10344], bl[10345], bl[10346], bl[10347], bl[10348], bl[10349], bl[10350], bl[10351], bl[10352], bl[10353], bl[10354], bl[10355], bl[10356], bl[10357], bl[10358], bl[10359], bl[10360], bl[10361], bl[10362], bl[10363], bl[10364], bl[10365], bl[10366], bl[10367], bl[10368], bl[10369], bl[10370], bl[10371], bl[10372], bl[10373], bl[10374], bl[10375], bl[10376], bl[10377], bl[10378], bl[10379], bl[10380], bl[10381], bl[10382], bl[10383], bl[10384], bl[10385], bl[10386], bl[10387], bl[10388], bl[10389], bl[10390], bl[10391], bl[10392], bl[10393], bl[10394], bl[10395], bl[10396], bl[10397], bl[10398], bl[10399], bl[10400], bl[10401], bl[10402], bl[10403], bl[10404], bl[10405], bl[10406], bl[10407], bl[10408], bl[10409], bl[10410], bl[10411], bl[10412], bl[10413], bl[10414], bl[10415], bl[10416], bl[10417], bl[10418], bl[10419], bl[10420], bl[10421], bl[10422], bl[10423], bl[11444], bl[11445], bl[11446], bl[11447], bl[11448], bl[11449], bl[11450], bl[11451], bl[11452], bl[11453], bl[11454], bl[11455], bl[11456], bl[11457], bl[11458], bl[11459], bl[11460], bl[11461], bl[11462], bl[11463], bl[11464], bl[11465], bl[11466], bl[11467], bl[11468], bl[11469], bl[11470], bl[11471], bl[11472], bl[11473], bl[11474], bl[11475], bl[11476], bl[11477], bl[11478], bl[11479], bl[11480], bl[11481], bl[11482], bl[11483], bl[11484], bl[11485], bl[11486], bl[11487], bl[11488], bl[11489], bl[11490], bl[11491], bl[11492], bl[11493], bl[11494], bl[11495], bl[11496], bl[11497], bl[11498], bl[11499], bl[11500], bl[11501], bl[11502], bl[11503], bl[11504], bl[11505], bl[11506], bl[11507], bl[11508], bl[11509], bl[11510], bl[11511], bl[11512], bl[11513], bl[11514], bl[11515], bl[11516], bl[11517], bl[11518], bl[11519], bl[11520], bl[11521], bl[11522], bl[11523]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    tile tile_2__4_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_0__3__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_0__3__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_0__3__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_1__2__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_1__2__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_1__2__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_0__2__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_0__2__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_0__2__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_0__2__grid_top_r_in[1]),
        .grid_left_in(grid_clb_1__3__grid_left_in),
        .grid_bottom_in(grid_clb_1__3__grid_bottom_in),
        .chanx_left_in(sb_0__1__2_chanx_right_out),
        .chanx_left_out(cbx_1__1__2_chanx_left_out),
        .grid_top_out(grid_clb_1__4__grid_bottom_in),
        .chany_bottom_in(sb_1__1__1_chany_top_out),
        .chany_bottom_out(cby_1__1__2_chany_bottom_out),
        .grid_right_out(grid_clb_2__3__grid_left_in),
        .chany_top_in_0(cby_1__1__3_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__5_chanx_left_out),
        .chany_top_out_0(sb_1__1__2_chany_top_out),
        .chanx_right_out_0(sb_1__1__2_chanx_right_out),
        .grid_top_r_in(sb_1__3__grid_top_r_in),
        .grid_top_l_in(sb_1__3__grid_top_l_in),
        .grid_right_t_in(sb_1__3__grid_right_t_in),
        .grid_right_b_in(sb_1__3__grid_right_b_in),
        .grid_bottom_r_in(sb_1__2__grid_top_r_in),
        .grid_bottom_l_in(sb_1__2__grid_top_l_in),
        .grid_left_t_in(sb_0__3__grid_right_t_in),
        .grid_left_b_in(sb_0__3__grid_right_b_in),
        .bl({bl[11684], bl[11685], bl[11686], bl[11687], bl[11688], bl[11689], bl[11690], bl[11691], bl[11692], bl[11693], bl[11694], bl[11695], bl[11696], bl[11697], bl[11698], bl[11699], bl[11700], bl[11701], bl[11702], bl[11703], bl[11704], bl[11705], bl[11706], bl[11707], bl[11708], bl[11709], bl[11710], bl[11711], bl[11712], bl[11713], bl[11714], bl[11715], bl[11716], bl[11717], bl[11718], bl[11719], bl[11720], bl[11721], bl[11722], bl[11723], bl[11724], bl[11725], bl[11726], bl[11727], bl[11728], bl[11729], bl[11730], bl[11731], bl[11732], bl[11733], bl[11734], bl[11735], bl[11736], bl[11737], bl[11738], bl[11739], bl[11740], bl[11741], bl[11742], bl[11743], bl[11744], bl[11745], bl[11746], bl[11747], bl[11748], bl[11749], bl[11750], bl[11751], bl[11752], bl[11753], bl[11754], bl[11755], bl[11756], bl[11757], bl[11758], bl[11759], bl[11760], bl[11761], bl[11762], bl[11763], bl[11764], bl[11765], bl[11766], bl[11767], bl[11768], bl[11769], bl[11770], bl[11771], bl[11772], bl[11773], bl[11774], bl[11775], bl[11776], bl[11777], bl[11778], bl[11779], bl[11780], bl[11781], bl[11782], bl[11783], bl[11784], bl[11785], bl[11786], bl[11787], bl[11788], bl[11789], bl[11790], bl[11791], bl[11792], bl[11793], bl[11794], bl[11795], bl[11796], bl[11797], bl[11798], bl[11799], bl[11800], bl[11801], bl[11802], bl[11803], bl[11804], bl[11805], bl[11806], bl[11807], bl[11808], bl[11809], bl[11810], bl[11811], bl[11812], bl[11813], bl[11814], bl[11815], bl[11816], bl[11817], bl[11818], bl[11819], bl[11820], bl[11821], bl[11822], bl[11823], bl[11824], bl[11825], bl[11826], bl[11827], bl[11828], bl[11829], bl[11830], bl[11831], bl[11832], bl[11833], bl[11834], bl[11835], bl[11836], bl[11837], bl[11838], bl[11839], bl[11840], bl[11841], bl[11842], bl[11843], bl[11844], bl[11845], bl[11846], bl[11847], bl[11848], bl[11849], bl[11850], bl[11851], bl[11852], bl[11853], bl[11854], bl[11855], bl[11856], bl[11857], bl[11858], bl[11859], bl[11860], bl[11861], bl[11862], bl[11863], bl[11864], bl[11865], bl[11866], bl[11867], bl[11868], bl[11869], bl[11870], bl[11871], bl[11872], bl[11873], bl[11874], bl[11875], bl[11876], bl[11877], bl[11878], bl[11879], bl[11880], bl[11881], bl[11882], bl[11883], bl[11884], bl[11885], bl[11886], bl[11887], bl[11888], bl[11889], bl[11890], bl[11891], bl[11892], bl[11893], bl[11894], bl[11895], bl[11896], bl[11897], bl[11898], bl[11899], bl[11900], bl[11901], bl[11902], bl[11903], bl[11904], bl[11905], bl[11906], bl[11907], bl[11908], bl[11909], bl[11910], bl[11911], bl[11912], bl[11913], bl[11914], bl[11915], bl[11916], bl[11917], bl[11918], bl[11919], bl[11920], bl[11921], bl[11922], bl[11923], bl[11924], bl[11925], bl[11926], bl[11927], bl[11928], bl[11929], bl[11930], bl[11931], bl[11932], bl[11933], bl[11934], bl[11935], bl[11936], bl[11937], bl[11938], bl[11939], bl[11940], bl[11941], bl[11942], bl[11943], bl[11944], bl[11945], bl[11946], bl[11947], bl[11948], bl[11949], bl[11950], bl[11951], bl[11952], bl[11953], bl[11954], bl[11955], bl[11956], bl[11957], bl[11958], bl[11959], bl[11960], bl[11961], bl[11962], bl[11963], bl[11964], bl[11965], bl[11966], bl[11967], bl[11968], bl[11969], bl[11970], bl[11971], bl[11972], bl[11973], bl[11974], bl[11975], bl[11976], bl[11977], bl[11978], bl[11979], bl[11980], bl[11981], bl[11982], bl[11983], bl[11984], bl[11985], bl[11986], bl[11987], bl[11988], bl[11989], bl[11990], bl[11991], bl[11992], bl[11993], bl[11994], bl[11995], bl[11996], bl[11997], bl[11998], bl[11999], bl[12000], bl[12001], bl[12002], bl[12003], bl[12004], bl[12005], bl[12006], bl[12007], bl[12008], bl[12009], bl[12010], bl[12011], bl[12012], bl[12013], bl[12014], bl[12015], bl[12016], bl[12017], bl[12018], bl[12019], bl[12020], bl[12021], bl[12022], bl[12023], bl[12024], bl[12025], bl[12026], bl[12027], bl[12028], bl[12029], bl[12030], bl[12031], bl[12032], bl[12033], bl[12034], bl[12035], bl[12036], bl[12037], bl[12038], bl[12039], bl[12040], bl[12041], bl[12042], bl[12043], bl[12044], bl[12045], bl[12046], bl[12047], bl[12048], bl[12049], bl[12050], bl[12051], bl[12052], bl[12053], bl[12054], bl[12055], bl[12056], bl[12057], bl[12058], bl[12059], bl[12060], bl[12061], bl[12062], bl[12063], bl[12064], bl[12065], bl[12066], bl[12067], bl[12068], bl[12069], bl[12070], bl[12071], bl[12072], bl[12073], bl[12074], bl[12075], bl[12076], bl[12077], bl[12078], bl[12079], bl[12080], bl[12081], bl[12082], bl[12083], bl[12084], bl[12085], bl[12086], bl[12087], bl[12088], bl[12089], bl[12090], bl[12091], bl[12092], bl[12093], bl[12094], bl[12095], bl[12096], bl[12097], bl[12098], bl[12099], bl[12100], bl[12101], bl[12102], bl[12103], bl[12104], bl[12105], bl[12106], bl[12107], bl[12108], bl[12109], bl[12110], bl[12111], bl[12112], bl[12113], bl[12114], bl[12115], bl[12116], bl[12117], bl[12118], bl[12119], bl[12120], bl[12121], bl[12122], bl[12123], bl[12124], bl[12125], bl[12126], bl[12127], bl[12128], bl[12129], bl[12130], bl[12131], bl[12132], bl[12133], bl[12134], bl[12135], bl[12136], bl[12137], bl[12138], bl[12139], bl[12140], bl[12141], bl[12142], bl[12143], bl[12144], bl[12145], bl[12146], bl[12147], bl[12148], bl[12149], bl[12150], bl[12151], bl[12152], bl[12153], bl[12154], bl[12155], bl[12156], bl[12157], bl[12158], bl[12159], bl[12160], bl[12161], bl[12162], bl[12163], bl[12164], bl[12165], bl[12166], bl[12167], bl[12168], bl[12169], bl[12170], bl[12171], bl[12172], bl[12173], bl[12174], bl[12175], bl[12176], bl[12177], bl[12178], bl[12179], bl[12180], bl[12181], bl[12182], bl[12183], bl[12184], bl[12185], bl[12186], bl[12187], bl[12188], bl[12189], bl[12190], bl[12191], bl[12192], bl[12193], bl[12194], bl[12195], bl[12196], bl[12197], bl[12198], bl[12199], bl[12200], bl[12201], bl[12202], bl[12203], bl[12204], bl[12205], bl[12206], bl[12207], bl[12208], bl[12209], bl[12210], bl[12211], bl[12212], bl[12213], bl[12214], bl[12215], bl[12216], bl[12217], bl[12218], bl[12219], bl[12220], bl[12221], bl[12222], bl[12223], bl[12224], bl[12225], bl[12226], bl[12227], bl[12228], bl[12229], bl[12230], bl[12231], bl[12232], bl[12233], bl[12234], bl[12235], bl[12236], bl[12237], bl[12238], bl[12239], bl[12240], bl[12241], bl[12242], bl[12243], bl[12244], bl[12245], bl[12246], bl[12247], bl[12248], bl[12249], bl[12250], bl[12251], bl[12252], bl[12253], bl[12254], bl[12255], bl[12256], bl[12257], bl[12258], bl[12259], bl[12260], bl[12261], bl[12262], bl[12263], bl[12264], bl[12265], bl[12266], bl[12267], bl[12268], bl[12269], bl[12270], bl[12271], bl[12272], bl[12273], bl[12274], bl[12275], bl[12276], bl[12277], bl[12278], bl[12279], bl[12280], bl[12281], bl[12282], bl[12283], bl[12284], bl[12285], bl[12286], bl[12287], bl[12288], bl[12289], bl[12290], bl[12291], bl[12292], bl[12293], bl[12294], bl[12295], bl[12296], bl[12297], bl[12298], bl[12299], bl[12300], bl[12301], bl[12302], bl[12303], bl[12304], bl[12305], bl[12306], bl[12307], bl[12308], bl[12309], bl[12310], bl[12311], bl[12312], bl[12313], bl[12314], bl[12315], bl[12316], bl[12317], bl[12318], bl[12319], bl[12320], bl[12321], bl[12322], bl[12323], bl[12324], bl[12325], bl[12326], bl[12327], bl[12328], bl[12329], bl[12330], bl[12331], bl[12332], bl[12333], bl[12334], bl[12335], bl[12336], bl[12337], bl[12338], bl[12339], bl[12340], bl[12341], bl[12342], bl[12343], bl[12344], bl[12345], bl[12346], bl[12347], bl[12348], bl[12349], bl[12350], bl[12351], bl[12352], bl[12353], bl[12354], bl[12355], bl[12356], bl[12357], bl[12358], bl[12359], bl[12360], bl[12361], bl[12362], bl[12363], bl[12364], bl[12365], bl[12366], bl[12367], bl[12368], bl[12369], bl[12370], bl[12371], bl[12372], bl[12373], bl[12374], bl[12375], bl[12376], bl[12377], bl[12378], bl[12379], bl[12380], bl[12381], bl[12382], bl[12383], bl[12384], bl[12385], bl[12386], bl[12387], bl[12388], bl[12389], bl[12390], bl[12391], bl[12392], bl[12393], bl[12394], bl[12395], bl[12396], bl[12397], bl[12398], bl[12399], bl[12400], bl[12401], bl[12402], bl[12403], bl[12404], bl[12405], bl[12406], bl[12407], bl[12408], bl[12409], bl[12410], bl[12411], bl[12412], bl[12413], bl[12414], bl[12415], bl[12416], bl[12417], bl[12418], bl[12419], bl[12420], bl[12421], bl[12422], bl[12423], bl[12424], bl[12425], bl[12426], bl[12427], bl[12428], bl[12429], bl[12430], bl[12431], bl[12432], bl[12433], bl[12434], bl[12435], bl[12436], bl[12437], bl[12438], bl[12439], bl[12440], bl[12441], bl[12442], bl[12443], bl[12444], bl[12445], bl[12446], bl[12447], bl[12448], bl[12449], bl[12450], bl[12451], bl[12452], bl[12453], bl[12454], bl[12455], bl[12456], bl[12457], bl[12458], bl[12459], bl[12460], bl[12461], bl[12462], bl[12463], bl[12464], bl[12465], bl[12466], bl[12467], bl[12468], bl[12469], bl[12470], bl[12471], bl[12472], bl[12473], bl[12474], bl[12475], bl[12476], bl[12477], bl[12478], bl[12479], bl[12480], bl[12481], bl[12482], bl[12483], bl[12484], bl[12485], bl[12486], bl[12487], bl[12488], bl[12489], bl[12490], bl[12491], bl[12492], bl[12493], bl[12494], bl[12495], bl[12496], bl[12497], bl[12498], bl[12499], bl[12500], bl[12501], bl[12502], bl[12503], bl[12504], bl[12505], bl[12506], bl[12507], bl[12508], bl[12509], bl[12510], bl[12511], bl[12512], bl[12513], bl[12514], bl[12515], bl[12516], bl[12517], bl[12518], bl[12519], bl[12520], bl[12521], bl[12522], bl[12523], bl[12524], bl[12525], bl[12526], bl[12527], bl[12528], bl[12529], bl[12530], bl[12531], bl[12532], bl[12533], bl[12534], bl[12535], bl[12536], bl[12537], bl[12538], bl[12539], bl[12540], bl[12541], bl[12542], bl[12543], bl[12544], bl[12545], bl[12546], bl[12547], bl[12548], bl[12549], bl[12550], bl[12551], bl[12552], bl[12553], bl[12554], bl[12555], bl[12556], bl[12557], bl[12558], bl[12559], bl[12560], bl[12561], bl[12562], bl[12563], bl[12564], bl[12565], bl[12566], bl[12567], bl[12568], bl[12569], bl[12570], bl[12571], bl[12572], bl[12573], bl[12574], bl[12575], bl[12576], bl[12577], bl[12578], bl[12579], bl[12580], bl[12581], bl[12582], bl[12583], bl[12584], bl[12585], bl[12586], bl[12587], bl[12588], bl[12589], bl[12590], bl[12591], bl[12592], bl[12593], bl[12594], bl[12595], bl[12596], bl[12597], bl[12598], bl[12599], bl[12600], bl[12601], bl[12602], bl[12603], bl[12604], bl[12605], bl[12606], bl[12607], bl[12608], bl[12609], bl[12610], bl[12611], bl[12612], bl[12613], bl[12614], bl[12615], bl[12616], bl[12617], bl[12618], bl[12619], bl[12620], bl[12621], bl[12622], bl[12623], bl[12624], bl[12625], bl[12626], bl[12627], bl[12628], bl[12629], bl[12630], bl[12631], bl[12632], bl[12633], bl[12634], bl[12635], bl[12636], bl[12637], bl[12638], bl[12639], bl[12640], bl[12641], bl[12642], bl[12643], bl[12644], bl[12645], bl[12646], bl[12647], bl[12648], bl[12649], bl[12650], bl[12651], bl[12652], bl[12653], bl[12654], bl[12655], bl[12656], bl[12657], bl[12658], bl[12659], bl[12660], bl[12661], bl[12662], bl[12663], bl[12664], bl[12665], bl[12666], bl[12667], bl[12668], bl[12669], bl[12670], bl[12671], bl[12672], bl[12673], bl[12674], bl[12675], bl[12676], bl[12677], bl[12678], bl[12679], bl[12680], bl[12681], bl[12682], bl[12683], bl[12684], bl[12685], bl[12686], bl[12687], bl[12688], bl[12689], bl[12690], bl[12691], bl[12692], bl[12693], bl[12694], bl[12695], bl[12696], bl[12697], bl[12698], bl[12699], bl[12700], bl[12701], bl[12702], bl[12703], bl[20328], bl[20329], bl[20330], bl[20331], bl[20332], bl[20333], bl[20334], bl[20335], bl[20336], bl[20337], bl[20338], bl[20339], bl[20340], bl[20341], bl[20342], bl[20343], bl[20344], bl[20345], bl[20346], bl[20347], bl[20348], bl[20349], bl[20350], bl[20351], bl[20352], bl[20353], bl[20354], bl[20355], bl[20356], bl[20357], bl[20358], bl[20359], bl[20360], bl[20361], bl[20362], bl[20363], bl[20364], bl[20365], bl[20366], bl[20367], bl[20368], bl[20369], bl[20370], bl[20371], bl[20372], bl[20373], bl[20374], bl[20375], bl[20376], bl[20377], bl[20378], bl[20379], bl[20380], bl[20381], bl[20382], bl[20383], bl[20384], bl[20385], bl[20386], bl[20387], bl[20388], bl[20389], bl[20390], bl[20391], bl[20392], bl[20393], bl[20394], bl[20395], bl[20396], bl[20397], bl[20398], bl[20399], bl[20400], bl[20401], bl[20402], bl[20403], bl[20404], bl[20405], bl[20406], bl[20407], bl[11604], bl[11605], bl[11606], bl[11607], bl[11608], bl[11609], bl[11610], bl[11611], bl[11612], bl[11613], bl[11614], bl[11615], bl[11616], bl[11617], bl[11618], bl[11619], bl[11620], bl[11621], bl[11622], bl[11623], bl[11624], bl[11625], bl[11626], bl[11627], bl[11628], bl[11629], bl[11630], bl[11631], bl[11632], bl[11633], bl[11634], bl[11635], bl[11636], bl[11637], bl[11638], bl[11639], bl[11640], bl[11641], bl[11642], bl[11643], bl[11644], bl[11645], bl[11646], bl[11647], bl[11648], bl[11649], bl[11650], bl[11651], bl[11652], bl[11653], bl[11654], bl[11655], bl[11656], bl[11657], bl[11658], bl[11659], bl[11660], bl[11661], bl[11662], bl[11663], bl[11664], bl[11665], bl[11666], bl[11667], bl[11668], bl[11669], bl[11670], bl[11671], bl[11672], bl[11673], bl[11674], bl[11675], bl[11676], bl[11677], bl[11678], bl[11679], bl[11680], bl[11681], bl[11682], bl[11683], bl[20248], bl[20249], bl[20250], bl[20251], bl[20252], bl[20253], bl[20254], bl[20255], bl[20256], bl[20257], bl[20258], bl[20259], bl[20260], bl[20261], bl[20262], bl[20263], bl[20264], bl[20265], bl[20266], bl[20267], bl[20268], bl[20269], bl[20270], bl[20271], bl[20272], bl[20273], bl[20274], bl[20275], bl[20276], bl[20277], bl[20278], bl[20279], bl[20280], bl[20281], bl[20282], bl[20283], bl[20284], bl[20285], bl[20286], bl[20287], bl[20288], bl[20289], bl[20290], bl[20291], bl[20292], bl[20293], bl[20294], bl[20295], bl[20296], bl[20297], bl[20298], bl[20299], bl[20300], bl[20301], bl[20302], bl[20303], bl[20304], bl[20305], bl[20306], bl[20307], bl[20308], bl[20309], bl[20310], bl[20311], bl[20312], bl[20313], bl[20314], bl[20315], bl[20316], bl[20317], bl[20318], bl[20319], bl[20320], bl[20321], bl[20322], bl[20323], bl[20324], bl[20325], bl[20326], bl[20327]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    tile tile_3__2_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_1__1__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_1__1__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_1__1__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_2__0__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_2__0__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_2__0__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_1__0__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_1__0__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_1__0__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_1__0__grid_top_r_in[1]),
        .grid_left_in(grid_clb_2__1__grid_left_in),
        .grid_bottom_in(grid_clb_2__1__grid_bottom_in),
        .chanx_left_in(sb_1__1__0_chanx_right_out),
        .chanx_left_out(cbx_1__1__3_chanx_left_out),
        .grid_top_out(grid_clb_2__2__grid_bottom_in),
        .chany_bottom_in(sb_1__0__1_chany_top_out),
        .chany_bottom_out(cby_1__1__4_chany_bottom_out),
        .grid_right_out(grid_clb_3__1__grid_left_in),
        .chany_top_in_0(cby_1__1__5_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__6_chanx_left_out),
        .chany_top_out_0(sb_1__1__3_chany_top_out),
        .chanx_right_out_0(sb_1__1__3_chanx_right_out),
        .grid_top_r_in(sb_2__1__grid_top_r_in),
        .grid_top_l_in(sb_2__1__grid_top_l_in),
        .grid_right_t_in(sb_2__1__grid_right_t_in),
        .grid_right_b_in(sb_2__1__grid_right_b_in),
        .grid_bottom_r_in(sb_2__0__grid_top_r_in),
        .grid_bottom_l_in(sb_2__0__grid_top_l_in),
        .grid_left_t_in(sb_1__1__grid_right_t_in),
        .grid_left_b_in(sb_1__1__grid_right_b_in),
        .bl({bl[2898], bl[2899], bl[2900], bl[2901], bl[2902], bl[2903], bl[2904], bl[2905], bl[2906], bl[2907], bl[2908], bl[2909], bl[2910], bl[2911], bl[2912], bl[2913], bl[2914], bl[2915], bl[2916], bl[2917], bl[2918], bl[2919], bl[2920], bl[2921], bl[2922], bl[2923], bl[2924], bl[2925], bl[2926], bl[2927], bl[2928], bl[2929], bl[2930], bl[2931], bl[2932], bl[2933], bl[2934], bl[2935], bl[2936], bl[2937], bl[2938], bl[2939], bl[2940], bl[2941], bl[2942], bl[2943], bl[2944], bl[2945], bl[2946], bl[2947], bl[2948], bl[2949], bl[2950], bl[2951], bl[2952], bl[2953], bl[2954], bl[2955], bl[2956], bl[2957], bl[2958], bl[2959], bl[2960], bl[2961], bl[2962], bl[2963], bl[2964], bl[2965], bl[2966], bl[2967], bl[2968], bl[2969], bl[2970], bl[2971], bl[2972], bl[2973], bl[2974], bl[2975], bl[2976], bl[2977], bl[2978], bl[2979], bl[2980], bl[2981], bl[2982], bl[2983], bl[2984], bl[2985], bl[2986], bl[2987], bl[2988], bl[2989], bl[2990], bl[2991], bl[2992], bl[2993], bl[2994], bl[2995], bl[2996], bl[2997], bl[2998], bl[2999], bl[3000], bl[3001], bl[3002], bl[3003], bl[3004], bl[3005], bl[3006], bl[3007], bl[3008], bl[3009], bl[3010], bl[3011], bl[3012], bl[3013], bl[3014], bl[3015], bl[3016], bl[3017], bl[3018], bl[3019], bl[3020], bl[3021], bl[3022], bl[3023], bl[3024], bl[3025], bl[3026], bl[3027], bl[3028], bl[3029], bl[3030], bl[3031], bl[3032], bl[3033], bl[3034], bl[3035], bl[3036], bl[3037], bl[3038], bl[3039], bl[3040], bl[3041], bl[3042], bl[3043], bl[3044], bl[3045], bl[3046], bl[3047], bl[3048], bl[3049], bl[3050], bl[3051], bl[3052], bl[3053], bl[3054], bl[3055], bl[3056], bl[3057], bl[3058], bl[3059], bl[3060], bl[3061], bl[3062], bl[3063], bl[3064], bl[3065], bl[3066], bl[3067], bl[3068], bl[3069], bl[3070], bl[3071], bl[3072], bl[3073], bl[3074], bl[3075], bl[3076], bl[3077], bl[3078], bl[3079], bl[3080], bl[3081], bl[3082], bl[3083], bl[3084], bl[3085], bl[3086], bl[3087], bl[3088], bl[3089], bl[3090], bl[3091], bl[3092], bl[3093], bl[3094], bl[3095], bl[3096], bl[3097], bl[3098], bl[3099], bl[3100], bl[3101], bl[3102], bl[3103], bl[3104], bl[3105], bl[3106], bl[3107], bl[3108], bl[3109], bl[3110], bl[3111], bl[3112], bl[3113], bl[3114], bl[3115], bl[3116], bl[3117], bl[3118], bl[3119], bl[3120], bl[3121], bl[3122], bl[3123], bl[3124], bl[3125], bl[3126], bl[3127], bl[3128], bl[3129], bl[3130], bl[3131], bl[3132], bl[3133], bl[3134], bl[3135], bl[3136], bl[3137], bl[3138], bl[3139], bl[3140], bl[3141], bl[3142], bl[3143], bl[3144], bl[3145], bl[3146], bl[3147], bl[3148], bl[3149], bl[3150], bl[3151], bl[3152], bl[3153], bl[3154], bl[3155], bl[3156], bl[3157], bl[3158], bl[3159], bl[3160], bl[3161], bl[3162], bl[3163], bl[3164], bl[3165], bl[3166], bl[3167], bl[3168], bl[3169], bl[3170], bl[3171], bl[3172], bl[3173], bl[3174], bl[3175], bl[3176], bl[3177], bl[3178], bl[3179], bl[3180], bl[3181], bl[3182], bl[3183], bl[3184], bl[3185], bl[3186], bl[3187], bl[3188], bl[3189], bl[3190], bl[3191], bl[3192], bl[3193], bl[3194], bl[3195], bl[3196], bl[3197], bl[3198], bl[3199], bl[3200], bl[3201], bl[3202], bl[3203], bl[3204], bl[3205], bl[3206], bl[3207], bl[3208], bl[3209], bl[3210], bl[3211], bl[3212], bl[3213], bl[3214], bl[3215], bl[3216], bl[3217], bl[3218], bl[3219], bl[3220], bl[3221], bl[3222], bl[3223], bl[3224], bl[3225], bl[3226], bl[3227], bl[3228], bl[3229], bl[3230], bl[3231], bl[3232], bl[3233], bl[3234], bl[3235], bl[3236], bl[3237], bl[3238], bl[3239], bl[3240], bl[3241], bl[3242], bl[3243], bl[3244], bl[3245], bl[3246], bl[3247], bl[3248], bl[3249], bl[3250], bl[3251], bl[3252], bl[3253], bl[3254], bl[3255], bl[3256], bl[3257], bl[3258], bl[3259], bl[3260], bl[3261], bl[3262], bl[3263], bl[3264], bl[3265], bl[3266], bl[3267], bl[3268], bl[3269], bl[3270], bl[3271], bl[3272], bl[3273], bl[3274], bl[3275], bl[3276], bl[3277], bl[3278], bl[3279], bl[3280], bl[3281], bl[3282], bl[3283], bl[3284], bl[3285], bl[3286], bl[3287], bl[3288], bl[3289], bl[3290], bl[3291], bl[3292], bl[3293], bl[3294], bl[3295], bl[3296], bl[3297], bl[3298], bl[3299], bl[3300], bl[3301], bl[3302], bl[3303], bl[3304], bl[3305], bl[3306], bl[3307], bl[3308], bl[3309], bl[3310], bl[3311], bl[3312], bl[3313], bl[3314], bl[3315], bl[3316], bl[3317], bl[3318], bl[3319], bl[3320], bl[3321], bl[3322], bl[3323], bl[3324], bl[3325], bl[3326], bl[3327], bl[3328], bl[3329], bl[3330], bl[3331], bl[3332], bl[3333], bl[3334], bl[3335], bl[3336], bl[3337], bl[3338], bl[3339], bl[3340], bl[3341], bl[3342], bl[3343], bl[3344], bl[3345], bl[3346], bl[3347], bl[3348], bl[3349], bl[3350], bl[3351], bl[3352], bl[3353], bl[3354], bl[3355], bl[3356], bl[3357], bl[3358], bl[3359], bl[3360], bl[3361], bl[3362], bl[3363], bl[3364], bl[3365], bl[3366], bl[3367], bl[3368], bl[3369], bl[3370], bl[3371], bl[3372], bl[3373], bl[3374], bl[3375], bl[3376], bl[3377], bl[3378], bl[3379], bl[3380], bl[3381], bl[3382], bl[3383], bl[3384], bl[3385], bl[3386], bl[3387], bl[3388], bl[3389], bl[3390], bl[3391], bl[3392], bl[3393], bl[3394], bl[3395], bl[3396], bl[3397], bl[3398], bl[3399], bl[3400], bl[3401], bl[3402], bl[3403], bl[3404], bl[3405], bl[3406], bl[3407], bl[3408], bl[3409], bl[3410], bl[3411], bl[3412], bl[3413], bl[3414], bl[3415], bl[3416], bl[3417], bl[3418], bl[3419], bl[3420], bl[3421], bl[3422], bl[3423], bl[3424], bl[3425], bl[3426], bl[3427], bl[3428], bl[3429], bl[3430], bl[3431], bl[3432], bl[3433], bl[3434], bl[3435], bl[3436], bl[3437], bl[3438], bl[3439], bl[3440], bl[3441], bl[3442], bl[3443], bl[3444], bl[3445], bl[3446], bl[3447], bl[3448], bl[3449], bl[3450], bl[3451], bl[3452], bl[3453], bl[3454], bl[3455], bl[3456], bl[3457], bl[3458], bl[3459], bl[3460], bl[3461], bl[3462], bl[3463], bl[3464], bl[3465], bl[3466], bl[3467], bl[3468], bl[3469], bl[3470], bl[3471], bl[3472], bl[3473], bl[3474], bl[3475], bl[3476], bl[3477], bl[3478], bl[3479], bl[3480], bl[3481], bl[3482], bl[3483], bl[3484], bl[3485], bl[3486], bl[3487], bl[3488], bl[3489], bl[3490], bl[3491], bl[3492], bl[3493], bl[3494], bl[3495], bl[3496], bl[3497], bl[3498], bl[3499], bl[3500], bl[3501], bl[3502], bl[3503], bl[3504], bl[3505], bl[3506], bl[3507], bl[3508], bl[3509], bl[3510], bl[3511], bl[3512], bl[3513], bl[3514], bl[3515], bl[3516], bl[3517], bl[3518], bl[3519], bl[3520], bl[3521], bl[3522], bl[3523], bl[3524], bl[3525], bl[3526], bl[3527], bl[3528], bl[3529], bl[3530], bl[3531], bl[3532], bl[3533], bl[3534], bl[3535], bl[3536], bl[3537], bl[3538], bl[3539], bl[3540], bl[3541], bl[3542], bl[3543], bl[3544], bl[3545], bl[3546], bl[3547], bl[3548], bl[3549], bl[3550], bl[3551], bl[3552], bl[3553], bl[3554], bl[3555], bl[3556], bl[3557], bl[3558], bl[3559], bl[3560], bl[3561], bl[3562], bl[3563], bl[3564], bl[3565], bl[3566], bl[3567], bl[3568], bl[3569], bl[3570], bl[3571], bl[3572], bl[3573], bl[3574], bl[3575], bl[3576], bl[3577], bl[3578], bl[3579], bl[3580], bl[3581], bl[3582], bl[3583], bl[3584], bl[3585], bl[3586], bl[3587], bl[3588], bl[3589], bl[3590], bl[3591], bl[3592], bl[3593], bl[3594], bl[3595], bl[3596], bl[3597], bl[3598], bl[3599], bl[3600], bl[3601], bl[3602], bl[3603], bl[3604], bl[3605], bl[3606], bl[3607], bl[3608], bl[3609], bl[3610], bl[3611], bl[3612], bl[3613], bl[3614], bl[3615], bl[3616], bl[3617], bl[3618], bl[3619], bl[3620], bl[3621], bl[3622], bl[3623], bl[3624], bl[3625], bl[3626], bl[3627], bl[3628], bl[3629], bl[3630], bl[3631], bl[3632], bl[3633], bl[3634], bl[3635], bl[3636], bl[3637], bl[3638], bl[3639], bl[3640], bl[3641], bl[3642], bl[3643], bl[3644], bl[3645], bl[3646], bl[3647], bl[3648], bl[3649], bl[3650], bl[3651], bl[3652], bl[3653], bl[3654], bl[3655], bl[3656], bl[3657], bl[3658], bl[3659], bl[3660], bl[3661], bl[3662], bl[3663], bl[3664], bl[3665], bl[3666], bl[3667], bl[3668], bl[3669], bl[3670], bl[3671], bl[3672], bl[3673], bl[3674], bl[3675], bl[3676], bl[3677], bl[3678], bl[3679], bl[3680], bl[3681], bl[3682], bl[3683], bl[3684], bl[3685], bl[3686], bl[3687], bl[3688], bl[3689], bl[3690], bl[3691], bl[3692], bl[3693], bl[3694], bl[3695], bl[3696], bl[3697], bl[3698], bl[3699], bl[3700], bl[3701], bl[3702], bl[3703], bl[3704], bl[3705], bl[3706], bl[3707], bl[3708], bl[3709], bl[3710], bl[3711], bl[3712], bl[3713], bl[3714], bl[3715], bl[3716], bl[3717], bl[3718], bl[3719], bl[3720], bl[3721], bl[3722], bl[3723], bl[3724], bl[3725], bl[3726], bl[3727], bl[3728], bl[3729], bl[3730], bl[3731], bl[3732], bl[3733], bl[3734], bl[3735], bl[3736], bl[3737], bl[3738], bl[3739], bl[3740], bl[3741], bl[3742], bl[3743], bl[3744], bl[3745], bl[3746], bl[3747], bl[3748], bl[3749], bl[3750], bl[3751], bl[3752], bl[3753], bl[3754], bl[3755], bl[3756], bl[3757], bl[3758], bl[3759], bl[3760], bl[3761], bl[3762], bl[3763], bl[3764], bl[3765], bl[3766], bl[3767], bl[3768], bl[3769], bl[3770], bl[3771], bl[3772], bl[3773], bl[3774], bl[3775], bl[3776], bl[3777], bl[3778], bl[3779], bl[3780], bl[3781], bl[3782], bl[3783], bl[3784], bl[3785], bl[3786], bl[3787], bl[3788], bl[3789], bl[3790], bl[3791], bl[3792], bl[3793], bl[3794], bl[3795], bl[3796], bl[3797], bl[3798], bl[3799], bl[3800], bl[3801], bl[3802], bl[3803], bl[3804], bl[3805], bl[3806], bl[3807], bl[3808], bl[3809], bl[3810], bl[3811], bl[3812], bl[3813], bl[3814], bl[3815], bl[3816], bl[3817], bl[3818], bl[3819], bl[3820], bl[3821], bl[3822], bl[3823], bl[3824], bl[3825], bl[3826], bl[3827], bl[3828], bl[3829], bl[3830], bl[3831], bl[3832], bl[3833], bl[3834], bl[3835], bl[3836], bl[3837], bl[3838], bl[3839], bl[3840], bl[3841], bl[3842], bl[3843], bl[3844], bl[3845], bl[3846], bl[3847], bl[3848], bl[3849], bl[3850], bl[3851], bl[3852], bl[3853], bl[3854], bl[3855], bl[3856], bl[3857], bl[3858], bl[3859], bl[3860], bl[3861], bl[3862], bl[3863], bl[3864], bl[3865], bl[3866], bl[3867], bl[3868], bl[3869], bl[3870], bl[3871], bl[3872], bl[3873], bl[3874], bl[3875], bl[3876], bl[3877], bl[3878], bl[3879], bl[3880], bl[3881], bl[3882], bl[3883], bl[3884], bl[3885], bl[3886], bl[3887], bl[3888], bl[3889], bl[3890], bl[3891], bl[3892], bl[3893], bl[3894], bl[3895], bl[3896], bl[3897], bl[3898], bl[3899], bl[3900], bl[3901], bl[3902], bl[3903], bl[3904], bl[3905], bl[3906], bl[3907], bl[3908], bl[3909], bl[3910], bl[3911], bl[3912], bl[3913], bl[3914], bl[3915], bl[3916], bl[3917], bl[9004], bl[9005], bl[9006], bl[9007], bl[9008], bl[9009], bl[9010], bl[9011], bl[9012], bl[9013], bl[9014], bl[9015], bl[9016], bl[9017], bl[9018], bl[9019], bl[9020], bl[9021], bl[9022], bl[9023], bl[9024], bl[9025], bl[9026], bl[9027], bl[9028], bl[9029], bl[9030], bl[9031], bl[9032], bl[9033], bl[9034], bl[9035], bl[9036], bl[9037], bl[9038], bl[9039], bl[9040], bl[9041], bl[9042], bl[9043], bl[9044], bl[9045], bl[9046], bl[9047], bl[9048], bl[9049], bl[9050], bl[9051], bl[9052], bl[9053], bl[9054], bl[9055], bl[9056], bl[9057], bl[9058], bl[9059], bl[9060], bl[9061], bl[9062], bl[9063], bl[9064], bl[9065], bl[9066], bl[9067], bl[9068], bl[9069], bl[9070], bl[9071], bl[9072], bl[9073], bl[9074], bl[9075], bl[9076], bl[9077], bl[9078], bl[9079], bl[9080], bl[9081], bl[9082], bl[9083], bl[2818], bl[2819], bl[2820], bl[2821], bl[2822], bl[2823], bl[2824], bl[2825], bl[2826], bl[2827], bl[2828], bl[2829], bl[2830], bl[2831], bl[2832], bl[2833], bl[2834], bl[2835], bl[2836], bl[2837], bl[2838], bl[2839], bl[2840], bl[2841], bl[2842], bl[2843], bl[2844], bl[2845], bl[2846], bl[2847], bl[2848], bl[2849], bl[2850], bl[2851], bl[2852], bl[2853], bl[2854], bl[2855], bl[2856], bl[2857], bl[2858], bl[2859], bl[2860], bl[2861], bl[2862], bl[2863], bl[2864], bl[2865], bl[2866], bl[2867], bl[2868], bl[2869], bl[2870], bl[2871], bl[2872], bl[2873], bl[2874], bl[2875], bl[2876], bl[2877], bl[2878], bl[2879], bl[2880], bl[2881], bl[2882], bl[2883], bl[2884], bl[2885], bl[2886], bl[2887], bl[2888], bl[2889], bl[2890], bl[2891], bl[2892], bl[2893], bl[2894], bl[2895], bl[2896], bl[2897], bl[8924], bl[8925], bl[8926], bl[8927], bl[8928], bl[8929], bl[8930], bl[8931], bl[8932], bl[8933], bl[8934], bl[8935], bl[8936], bl[8937], bl[8938], bl[8939], bl[8940], bl[8941], bl[8942], bl[8943], bl[8944], bl[8945], bl[8946], bl[8947], bl[8948], bl[8949], bl[8950], bl[8951], bl[8952], bl[8953], bl[8954], bl[8955], bl[8956], bl[8957], bl[8958], bl[8959], bl[8960], bl[8961], bl[8962], bl[8963], bl[8964], bl[8965], bl[8966], bl[8967], bl[8968], bl[8969], bl[8970], bl[8971], bl[8972], bl[8973], bl[8974], bl[8975], bl[8976], bl[8977], bl[8978], bl[8979], bl[8980], bl[8981], bl[8982], bl[8983], bl[8984], bl[8985], bl[8986], bl[8987], bl[8988], bl[8989], bl[8990], bl[8991], bl[8992], bl[8993], bl[8994], bl[8995], bl[8996], bl[8997], bl[8998], bl[8999], bl[9000], bl[9001], bl[9002], bl[9003]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    tile tile_3__3_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_1__2__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_1__2__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_1__2__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_2__1__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_2__1__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_2__1__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_1__1__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_1__1__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_1__1__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_1__1__grid_top_r_in[1]),
        .grid_left_in(grid_clb_2__2__grid_left_in),
        .grid_bottom_in(grid_clb_2__2__grid_bottom_in),
        .chanx_left_in(sb_1__1__1_chanx_right_out),
        .chanx_left_out(cbx_1__1__4_chanx_left_out),
        .grid_top_out(grid_clb_2__3__grid_bottom_in),
        .chany_bottom_in(sb_1__1__3_chany_top_out),
        .chany_bottom_out(cby_1__1__5_chany_bottom_out),
        .grid_right_out(grid_clb_3__2__grid_left_in),
        .chany_top_in_0(cby_1__1__6_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__7_chanx_left_out),
        .chany_top_out_0(sb_1__1__4_chany_top_out),
        .chanx_right_out_0(sb_1__1__4_chanx_right_out),
        .grid_top_r_in(sb_2__2__grid_top_r_in),
        .grid_top_l_in(sb_2__2__grid_top_l_in),
        .grid_right_t_in(sb_2__2__grid_right_t_in),
        .grid_right_b_in(sb_2__2__grid_right_b_in),
        .grid_bottom_r_in(sb_2__1__grid_top_r_in),
        .grid_bottom_l_in(sb_2__1__grid_top_l_in),
        .grid_left_t_in(sb_1__2__grid_right_t_in),
        .grid_left_b_in(sb_1__2__grid_right_b_in),
        .bl({bl[9164], bl[9165], bl[9166], bl[9167], bl[9168], bl[9169], bl[9170], bl[9171], bl[9172], bl[9173], bl[9174], bl[9175], bl[9176], bl[9177], bl[9178], bl[9179], bl[9180], bl[9181], bl[9182], bl[9183], bl[9184], bl[9185], bl[9186], bl[9187], bl[9188], bl[9189], bl[9190], bl[9191], bl[9192], bl[9193], bl[9194], bl[9195], bl[9196], bl[9197], bl[9198], bl[9199], bl[9200], bl[9201], bl[9202], bl[9203], bl[9204], bl[9205], bl[9206], bl[9207], bl[9208], bl[9209], bl[9210], bl[9211], bl[9212], bl[9213], bl[9214], bl[9215], bl[9216], bl[9217], bl[9218], bl[9219], bl[9220], bl[9221], bl[9222], bl[9223], bl[9224], bl[9225], bl[9226], bl[9227], bl[9228], bl[9229], bl[9230], bl[9231], bl[9232], bl[9233], bl[9234], bl[9235], bl[9236], bl[9237], bl[9238], bl[9239], bl[9240], bl[9241], bl[9242], bl[9243], bl[9244], bl[9245], bl[9246], bl[9247], bl[9248], bl[9249], bl[9250], bl[9251], bl[9252], bl[9253], bl[9254], bl[9255], bl[9256], bl[9257], bl[9258], bl[9259], bl[9260], bl[9261], bl[9262], bl[9263], bl[9264], bl[9265], bl[9266], bl[9267], bl[9268], bl[9269], bl[9270], bl[9271], bl[9272], bl[9273], bl[9274], bl[9275], bl[9276], bl[9277], bl[9278], bl[9279], bl[9280], bl[9281], bl[9282], bl[9283], bl[9284], bl[9285], bl[9286], bl[9287], bl[9288], bl[9289], bl[9290], bl[9291], bl[9292], bl[9293], bl[9294], bl[9295], bl[9296], bl[9297], bl[9298], bl[9299], bl[9300], bl[9301], bl[9302], bl[9303], bl[9304], bl[9305], bl[9306], bl[9307], bl[9308], bl[9309], bl[9310], bl[9311], bl[9312], bl[9313], bl[9314], bl[9315], bl[9316], bl[9317], bl[9318], bl[9319], bl[9320], bl[9321], bl[9322], bl[9323], bl[9324], bl[9325], bl[9326], bl[9327], bl[9328], bl[9329], bl[9330], bl[9331], bl[9332], bl[9333], bl[9334], bl[9335], bl[9336], bl[9337], bl[9338], bl[9339], bl[9340], bl[9341], bl[9342], bl[9343], bl[9344], bl[9345], bl[9346], bl[9347], bl[9348], bl[9349], bl[9350], bl[9351], bl[9352], bl[9353], bl[9354], bl[9355], bl[9356], bl[9357], bl[9358], bl[9359], bl[9360], bl[9361], bl[9362], bl[9363], bl[9364], bl[9365], bl[9366], bl[9367], bl[9368], bl[9369], bl[9370], bl[9371], bl[9372], bl[9373], bl[9374], bl[9375], bl[9376], bl[9377], bl[9378], bl[9379], bl[9380], bl[9381], bl[9382], bl[9383], bl[9384], bl[9385], bl[9386], bl[9387], bl[9388], bl[9389], bl[9390], bl[9391], bl[9392], bl[9393], bl[9394], bl[9395], bl[9396], bl[9397], bl[9398], bl[9399], bl[9400], bl[9401], bl[9402], bl[9403], bl[9404], bl[9405], bl[9406], bl[9407], bl[9408], bl[9409], bl[9410], bl[9411], bl[9412], bl[9413], bl[9414], bl[9415], bl[9416], bl[9417], bl[9418], bl[9419], bl[9420], bl[9421], bl[9422], bl[9423], bl[9424], bl[9425], bl[9426], bl[9427], bl[9428], bl[9429], bl[9430], bl[9431], bl[9432], bl[9433], bl[9434], bl[9435], bl[9436], bl[9437], bl[9438], bl[9439], bl[9440], bl[9441], bl[9442], bl[9443], bl[9444], bl[9445], bl[9446], bl[9447], bl[9448], bl[9449], bl[9450], bl[9451], bl[9452], bl[9453], bl[9454], bl[9455], bl[9456], bl[9457], bl[9458], bl[9459], bl[9460], bl[9461], bl[9462], bl[9463], bl[9464], bl[9465], bl[9466], bl[9467], bl[9468], bl[9469], bl[9470], bl[9471], bl[9472], bl[9473], bl[9474], bl[9475], bl[9476], bl[9477], bl[9478], bl[9479], bl[9480], bl[9481], bl[9482], bl[9483], bl[9484], bl[9485], bl[9486], bl[9487], bl[9488], bl[9489], bl[9490], bl[9491], bl[9492], bl[9493], bl[9494], bl[9495], bl[9496], bl[9497], bl[9498], bl[9499], bl[9500], bl[9501], bl[9502], bl[9503], bl[9504], bl[9505], bl[9506], bl[9507], bl[9508], bl[9509], bl[9510], bl[9511], bl[9512], bl[9513], bl[9514], bl[9515], bl[9516], bl[9517], bl[9518], bl[9519], bl[9520], bl[9521], bl[9522], bl[9523], bl[9524], bl[9525], bl[9526], bl[9527], bl[9528], bl[9529], bl[9530], bl[9531], bl[9532], bl[9533], bl[9534], bl[9535], bl[9536], bl[9537], bl[9538], bl[9539], bl[9540], bl[9541], bl[9542], bl[9543], bl[9544], bl[9545], bl[9546], bl[9547], bl[9548], bl[9549], bl[9550], bl[9551], bl[9552], bl[9553], bl[9554], bl[9555], bl[9556], bl[9557], bl[9558], bl[9559], bl[9560], bl[9561], bl[9562], bl[9563], bl[9564], bl[9565], bl[9566], bl[9567], bl[9568], bl[9569], bl[9570], bl[9571], bl[9572], bl[9573], bl[9574], bl[9575], bl[9576], bl[9577], bl[9578], bl[9579], bl[9580], bl[9581], bl[9582], bl[9583], bl[9584], bl[9585], bl[9586], bl[9587], bl[9588], bl[9589], bl[9590], bl[9591], bl[9592], bl[9593], bl[9594], bl[9595], bl[9596], bl[9597], bl[9598], bl[9599], bl[9600], bl[9601], bl[9602], bl[9603], bl[9604], bl[9605], bl[9606], bl[9607], bl[9608], bl[9609], bl[9610], bl[9611], bl[9612], bl[9613], bl[9614], bl[9615], bl[9616], bl[9617], bl[9618], bl[9619], bl[9620], bl[9621], bl[9622], bl[9623], bl[9624], bl[9625], bl[9626], bl[9627], bl[9628], bl[9629], bl[9630], bl[9631], bl[9632], bl[9633], bl[9634], bl[9635], bl[9636], bl[9637], bl[9638], bl[9639], bl[9640], bl[9641], bl[9642], bl[9643], bl[9644], bl[9645], bl[9646], bl[9647], bl[9648], bl[9649], bl[9650], bl[9651], bl[9652], bl[9653], bl[9654], bl[9655], bl[9656], bl[9657], bl[9658], bl[9659], bl[9660], bl[9661], bl[9662], bl[9663], bl[9664], bl[9665], bl[9666], bl[9667], bl[9668], bl[9669], bl[9670], bl[9671], bl[9672], bl[9673], bl[9674], bl[9675], bl[9676], bl[9677], bl[9678], bl[9679], bl[9680], bl[9681], bl[9682], bl[9683], bl[9684], bl[9685], bl[9686], bl[9687], bl[9688], bl[9689], bl[9690], bl[9691], bl[9692], bl[9693], bl[9694], bl[9695], bl[9696], bl[9697], bl[9698], bl[9699], bl[9700], bl[9701], bl[9702], bl[9703], bl[9704], bl[9705], bl[9706], bl[9707], bl[9708], bl[9709], bl[9710], bl[9711], bl[9712], bl[9713], bl[9714], bl[9715], bl[9716], bl[9717], bl[9718], bl[9719], bl[9720], bl[9721], bl[9722], bl[9723], bl[9724], bl[9725], bl[9726], bl[9727], bl[9728], bl[9729], bl[9730], bl[9731], bl[9732], bl[9733], bl[9734], bl[9735], bl[9736], bl[9737], bl[9738], bl[9739], bl[9740], bl[9741], bl[9742], bl[9743], bl[9744], bl[9745], bl[9746], bl[9747], bl[9748], bl[9749], bl[9750], bl[9751], bl[9752], bl[9753], bl[9754], bl[9755], bl[9756], bl[9757], bl[9758], bl[9759], bl[9760], bl[9761], bl[9762], bl[9763], bl[9764], bl[9765], bl[9766], bl[9767], bl[9768], bl[9769], bl[9770], bl[9771], bl[9772], bl[9773], bl[9774], bl[9775], bl[9776], bl[9777], bl[9778], bl[9779], bl[9780], bl[9781], bl[9782], bl[9783], bl[9784], bl[9785], bl[9786], bl[9787], bl[9788], bl[9789], bl[9790], bl[9791], bl[9792], bl[9793], bl[9794], bl[9795], bl[9796], bl[9797], bl[9798], bl[9799], bl[9800], bl[9801], bl[9802], bl[9803], bl[9804], bl[9805], bl[9806], bl[9807], bl[9808], bl[9809], bl[9810], bl[9811], bl[9812], bl[9813], bl[9814], bl[9815], bl[9816], bl[9817], bl[9818], bl[9819], bl[9820], bl[9821], bl[9822], bl[9823], bl[9824], bl[9825], bl[9826], bl[9827], bl[9828], bl[9829], bl[9830], bl[9831], bl[9832], bl[9833], bl[9834], bl[9835], bl[9836], bl[9837], bl[9838], bl[9839], bl[9840], bl[9841], bl[9842], bl[9843], bl[9844], bl[9845], bl[9846], bl[9847], bl[9848], bl[9849], bl[9850], bl[9851], bl[9852], bl[9853], bl[9854], bl[9855], bl[9856], bl[9857], bl[9858], bl[9859], bl[9860], bl[9861], bl[9862], bl[9863], bl[9864], bl[9865], bl[9866], bl[9867], bl[9868], bl[9869], bl[9870], bl[9871], bl[9872], bl[9873], bl[9874], bl[9875], bl[9876], bl[9877], bl[9878], bl[9879], bl[9880], bl[9881], bl[9882], bl[9883], bl[9884], bl[9885], bl[9886], bl[9887], bl[9888], bl[9889], bl[9890], bl[9891], bl[9892], bl[9893], bl[9894], bl[9895], bl[9896], bl[9897], bl[9898], bl[9899], bl[9900], bl[9901], bl[9902], bl[9903], bl[9904], bl[9905], bl[9906], bl[9907], bl[9908], bl[9909], bl[9910], bl[9911], bl[9912], bl[9913], bl[9914], bl[9915], bl[9916], bl[9917], bl[9918], bl[9919], bl[9920], bl[9921], bl[9922], bl[9923], bl[9924], bl[9925], bl[9926], bl[9927], bl[9928], bl[9929], bl[9930], bl[9931], bl[9932], bl[9933], bl[9934], bl[9935], bl[9936], bl[9937], bl[9938], bl[9939], bl[9940], bl[9941], bl[9942], bl[9943], bl[9944], bl[9945], bl[9946], bl[9947], bl[9948], bl[9949], bl[9950], bl[9951], bl[9952], bl[9953], bl[9954], bl[9955], bl[9956], bl[9957], bl[9958], bl[9959], bl[9960], bl[9961], bl[9962], bl[9963], bl[9964], bl[9965], bl[9966], bl[9967], bl[9968], bl[9969], bl[9970], bl[9971], bl[9972], bl[9973], bl[9974], bl[9975], bl[9976], bl[9977], bl[9978], bl[9979], bl[9980], bl[9981], bl[9982], bl[9983], bl[9984], bl[9985], bl[9986], bl[9987], bl[9988], bl[9989], bl[9990], bl[9991], bl[9992], bl[9993], bl[9994], bl[9995], bl[9996], bl[9997], bl[9998], bl[9999], bl[10000], bl[10001], bl[10002], bl[10003], bl[10004], bl[10005], bl[10006], bl[10007], bl[10008], bl[10009], bl[10010], bl[10011], bl[10012], bl[10013], bl[10014], bl[10015], bl[10016], bl[10017], bl[10018], bl[10019], bl[10020], bl[10021], bl[10022], bl[10023], bl[10024], bl[10025], bl[10026], bl[10027], bl[10028], bl[10029], bl[10030], bl[10031], bl[10032], bl[10033], bl[10034], bl[10035], bl[10036], bl[10037], bl[10038], bl[10039], bl[10040], bl[10041], bl[10042], bl[10043], bl[10044], bl[10045], bl[10046], bl[10047], bl[10048], bl[10049], bl[10050], bl[10051], bl[10052], bl[10053], bl[10054], bl[10055], bl[10056], bl[10057], bl[10058], bl[10059], bl[10060], bl[10061], bl[10062], bl[10063], bl[10064], bl[10065], bl[10066], bl[10067], bl[10068], bl[10069], bl[10070], bl[10071], bl[10072], bl[10073], bl[10074], bl[10075], bl[10076], bl[10077], bl[10078], bl[10079], bl[10080], bl[10081], bl[10082], bl[10083], bl[10084], bl[10085], bl[10086], bl[10087], bl[10088], bl[10089], bl[10090], bl[10091], bl[10092], bl[10093], bl[10094], bl[10095], bl[10096], bl[10097], bl[10098], bl[10099], bl[10100], bl[10101], bl[10102], bl[10103], bl[10104], bl[10105], bl[10106], bl[10107], bl[10108], bl[10109], bl[10110], bl[10111], bl[10112], bl[10113], bl[10114], bl[10115], bl[10116], bl[10117], bl[10118], bl[10119], bl[10120], bl[10121], bl[10122], bl[10123], bl[10124], bl[10125], bl[10126], bl[10127], bl[10128], bl[10129], bl[10130], bl[10131], bl[10132], bl[10133], bl[10134], bl[10135], bl[10136], bl[10137], bl[10138], bl[10139], bl[10140], bl[10141], bl[10142], bl[10143], bl[10144], bl[10145], bl[10146], bl[10147], bl[10148], bl[10149], bl[10150], bl[10151], bl[10152], bl[10153], bl[10154], bl[10155], bl[10156], bl[10157], bl[10158], bl[10159], bl[10160], bl[10161], bl[10162], bl[10163], bl[10164], bl[10165], bl[10166], bl[10167], bl[10168], bl[10169], bl[10170], bl[10171], bl[10172], bl[10173], bl[10174], bl[10175], bl[10176], bl[10177], bl[10178], bl[10179], bl[10180], bl[10181], bl[10182], bl[10183], bl[12784], bl[12785], bl[12786], bl[12787], bl[12788], bl[12789], bl[12790], bl[12791], bl[12792], bl[12793], bl[12794], bl[12795], bl[12796], bl[12797], bl[12798], bl[12799], bl[12800], bl[12801], bl[12802], bl[12803], bl[12804], bl[12805], bl[12806], bl[12807], bl[12808], bl[12809], bl[12810], bl[12811], bl[12812], bl[12813], bl[12814], bl[12815], bl[12816], bl[12817], bl[12818], bl[12819], bl[12820], bl[12821], bl[12822], bl[12823], bl[12824], bl[12825], bl[12826], bl[12827], bl[12828], bl[12829], bl[12830], bl[12831], bl[12832], bl[12833], bl[12834], bl[12835], bl[12836], bl[12837], bl[12838], bl[12839], bl[12840], bl[12841], bl[12842], bl[12843], bl[12844], bl[12845], bl[12846], bl[12847], bl[12848], bl[12849], bl[12850], bl[12851], bl[12852], bl[12853], bl[12854], bl[12855], bl[12856], bl[12857], bl[12858], bl[12859], bl[12860], bl[12861], bl[12862], bl[12863], bl[9084], bl[9085], bl[9086], bl[9087], bl[9088], bl[9089], bl[9090], bl[9091], bl[9092], bl[9093], bl[9094], bl[9095], bl[9096], bl[9097], bl[9098], bl[9099], bl[9100], bl[9101], bl[9102], bl[9103], bl[9104], bl[9105], bl[9106], bl[9107], bl[9108], bl[9109], bl[9110], bl[9111], bl[9112], bl[9113], bl[9114], bl[9115], bl[9116], bl[9117], bl[9118], bl[9119], bl[9120], bl[9121], bl[9122], bl[9123], bl[9124], bl[9125], bl[9126], bl[9127], bl[9128], bl[9129], bl[9130], bl[9131], bl[9132], bl[9133], bl[9134], bl[9135], bl[9136], bl[9137], bl[9138], bl[9139], bl[9140], bl[9141], bl[9142], bl[9143], bl[9144], bl[9145], bl[9146], bl[9147], bl[9148], bl[9149], bl[9150], bl[9151], bl[9152], bl[9153], bl[9154], bl[9155], bl[9156], bl[9157], bl[9158], bl[9159], bl[9160], bl[9161], bl[9162], bl[9163], bl[12704], bl[12705], bl[12706], bl[12707], bl[12708], bl[12709], bl[12710], bl[12711], bl[12712], bl[12713], bl[12714], bl[12715], bl[12716], bl[12717], bl[12718], bl[12719], bl[12720], bl[12721], bl[12722], bl[12723], bl[12724], bl[12725], bl[12726], bl[12727], bl[12728], bl[12729], bl[12730], bl[12731], bl[12732], bl[12733], bl[12734], bl[12735], bl[12736], bl[12737], bl[12738], bl[12739], bl[12740], bl[12741], bl[12742], bl[12743], bl[12744], bl[12745], bl[12746], bl[12747], bl[12748], bl[12749], bl[12750], bl[12751], bl[12752], bl[12753], bl[12754], bl[12755], bl[12756], bl[12757], bl[12758], bl[12759], bl[12760], bl[12761], bl[12762], bl[12763], bl[12764], bl[12765], bl[12766], bl[12767], bl[12768], bl[12769], bl[12770], bl[12771], bl[12772], bl[12773], bl[12774], bl[12775], bl[12776], bl[12777], bl[12778], bl[12779], bl[12780], bl[12781], bl[12782], bl[12783]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    tile tile_3__4_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_1__3__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_1__3__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_1__3__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_2__2__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_2__2__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_2__2__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_1__2__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_1__2__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_1__2__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_1__2__grid_top_r_in[1]),
        .grid_left_in(grid_clb_2__3__grid_left_in),
        .grid_bottom_in(grid_clb_2__3__grid_bottom_in),
        .chanx_left_in(sb_1__1__2_chanx_right_out),
        .chanx_left_out(cbx_1__1__5_chanx_left_out),
        .grid_top_out(grid_clb_2__4__grid_bottom_in),
        .chany_bottom_in(sb_1__1__4_chany_top_out),
        .chany_bottom_out(cby_1__1__6_chany_bottom_out),
        .grid_right_out(grid_clb_3__3__grid_left_in),
        .chany_top_in_0(cby_1__1__7_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__8_chanx_left_out),
        .chany_top_out_0(sb_1__1__5_chany_top_out),
        .chanx_right_out_0(sb_1__1__5_chanx_right_out),
        .grid_top_r_in(sb_2__3__grid_top_r_in),
        .grid_top_l_in(sb_2__3__grid_top_l_in),
        .grid_right_t_in(sb_2__3__grid_right_t_in),
        .grid_right_b_in(sb_2__3__grid_right_b_in),
        .grid_bottom_r_in(sb_2__2__grid_top_r_in),
        .grid_bottom_l_in(sb_2__2__grid_top_l_in),
        .grid_left_t_in(sb_1__3__grid_right_t_in),
        .grid_left_b_in(sb_1__3__grid_right_b_in),
        .bl({bl[12944], bl[12945], bl[12946], bl[12947], bl[12948], bl[12949], bl[12950], bl[12951], bl[12952], bl[12953], bl[12954], bl[12955], bl[12956], bl[12957], bl[12958], bl[12959], bl[12960], bl[12961], bl[12962], bl[12963], bl[12964], bl[12965], bl[12966], bl[12967], bl[12968], bl[12969], bl[12970], bl[12971], bl[12972], bl[12973], bl[12974], bl[12975], bl[12976], bl[12977], bl[12978], bl[12979], bl[12980], bl[12981], bl[12982], bl[12983], bl[12984], bl[12985], bl[12986], bl[12987], bl[12988], bl[12989], bl[12990], bl[12991], bl[12992], bl[12993], bl[12994], bl[12995], bl[12996], bl[12997], bl[12998], bl[12999], bl[13000], bl[13001], bl[13002], bl[13003], bl[13004], bl[13005], bl[13006], bl[13007], bl[13008], bl[13009], bl[13010], bl[13011], bl[13012], bl[13013], bl[13014], bl[13015], bl[13016], bl[13017], bl[13018], bl[13019], bl[13020], bl[13021], bl[13022], bl[13023], bl[13024], bl[13025], bl[13026], bl[13027], bl[13028], bl[13029], bl[13030], bl[13031], bl[13032], bl[13033], bl[13034], bl[13035], bl[13036], bl[13037], bl[13038], bl[13039], bl[13040], bl[13041], bl[13042], bl[13043], bl[13044], bl[13045], bl[13046], bl[13047], bl[13048], bl[13049], bl[13050], bl[13051], bl[13052], bl[13053], bl[13054], bl[13055], bl[13056], bl[13057], bl[13058], bl[13059], bl[13060], bl[13061], bl[13062], bl[13063], bl[13064], bl[13065], bl[13066], bl[13067], bl[13068], bl[13069], bl[13070], bl[13071], bl[13072], bl[13073], bl[13074], bl[13075], bl[13076], bl[13077], bl[13078], bl[13079], bl[13080], bl[13081], bl[13082], bl[13083], bl[13084], bl[13085], bl[13086], bl[13087], bl[13088], bl[13089], bl[13090], bl[13091], bl[13092], bl[13093], bl[13094], bl[13095], bl[13096], bl[13097], bl[13098], bl[13099], bl[13100], bl[13101], bl[13102], bl[13103], bl[13104], bl[13105], bl[13106], bl[13107], bl[13108], bl[13109], bl[13110], bl[13111], bl[13112], bl[13113], bl[13114], bl[13115], bl[13116], bl[13117], bl[13118], bl[13119], bl[13120], bl[13121], bl[13122], bl[13123], bl[13124], bl[13125], bl[13126], bl[13127], bl[13128], bl[13129], bl[13130], bl[13131], bl[13132], bl[13133], bl[13134], bl[13135], bl[13136], bl[13137], bl[13138], bl[13139], bl[13140], bl[13141], bl[13142], bl[13143], bl[13144], bl[13145], bl[13146], bl[13147], bl[13148], bl[13149], bl[13150], bl[13151], bl[13152], bl[13153], bl[13154], bl[13155], bl[13156], bl[13157], bl[13158], bl[13159], bl[13160], bl[13161], bl[13162], bl[13163], bl[13164], bl[13165], bl[13166], bl[13167], bl[13168], bl[13169], bl[13170], bl[13171], bl[13172], bl[13173], bl[13174], bl[13175], bl[13176], bl[13177], bl[13178], bl[13179], bl[13180], bl[13181], bl[13182], bl[13183], bl[13184], bl[13185], bl[13186], bl[13187], bl[13188], bl[13189], bl[13190], bl[13191], bl[13192], bl[13193], bl[13194], bl[13195], bl[13196], bl[13197], bl[13198], bl[13199], bl[13200], bl[13201], bl[13202], bl[13203], bl[13204], bl[13205], bl[13206], bl[13207], bl[13208], bl[13209], bl[13210], bl[13211], bl[13212], bl[13213], bl[13214], bl[13215], bl[13216], bl[13217], bl[13218], bl[13219], bl[13220], bl[13221], bl[13222], bl[13223], bl[13224], bl[13225], bl[13226], bl[13227], bl[13228], bl[13229], bl[13230], bl[13231], bl[13232], bl[13233], bl[13234], bl[13235], bl[13236], bl[13237], bl[13238], bl[13239], bl[13240], bl[13241], bl[13242], bl[13243], bl[13244], bl[13245], bl[13246], bl[13247], bl[13248], bl[13249], bl[13250], bl[13251], bl[13252], bl[13253], bl[13254], bl[13255], bl[13256], bl[13257], bl[13258], bl[13259], bl[13260], bl[13261], bl[13262], bl[13263], bl[13264], bl[13265], bl[13266], bl[13267], bl[13268], bl[13269], bl[13270], bl[13271], bl[13272], bl[13273], bl[13274], bl[13275], bl[13276], bl[13277], bl[13278], bl[13279], bl[13280], bl[13281], bl[13282], bl[13283], bl[13284], bl[13285], bl[13286], bl[13287], bl[13288], bl[13289], bl[13290], bl[13291], bl[13292], bl[13293], bl[13294], bl[13295], bl[13296], bl[13297], bl[13298], bl[13299], bl[13300], bl[13301], bl[13302], bl[13303], bl[13304], bl[13305], bl[13306], bl[13307], bl[13308], bl[13309], bl[13310], bl[13311], bl[13312], bl[13313], bl[13314], bl[13315], bl[13316], bl[13317], bl[13318], bl[13319], bl[13320], bl[13321], bl[13322], bl[13323], bl[13324], bl[13325], bl[13326], bl[13327], bl[13328], bl[13329], bl[13330], bl[13331], bl[13332], bl[13333], bl[13334], bl[13335], bl[13336], bl[13337], bl[13338], bl[13339], bl[13340], bl[13341], bl[13342], bl[13343], bl[13344], bl[13345], bl[13346], bl[13347], bl[13348], bl[13349], bl[13350], bl[13351], bl[13352], bl[13353], bl[13354], bl[13355], bl[13356], bl[13357], bl[13358], bl[13359], bl[13360], bl[13361], bl[13362], bl[13363], bl[13364], bl[13365], bl[13366], bl[13367], bl[13368], bl[13369], bl[13370], bl[13371], bl[13372], bl[13373], bl[13374], bl[13375], bl[13376], bl[13377], bl[13378], bl[13379], bl[13380], bl[13381], bl[13382], bl[13383], bl[13384], bl[13385], bl[13386], bl[13387], bl[13388], bl[13389], bl[13390], bl[13391], bl[13392], bl[13393], bl[13394], bl[13395], bl[13396], bl[13397], bl[13398], bl[13399], bl[13400], bl[13401], bl[13402], bl[13403], bl[13404], bl[13405], bl[13406], bl[13407], bl[13408], bl[13409], bl[13410], bl[13411], bl[13412], bl[13413], bl[13414], bl[13415], bl[13416], bl[13417], bl[13418], bl[13419], bl[13420], bl[13421], bl[13422], bl[13423], bl[13424], bl[13425], bl[13426], bl[13427], bl[13428], bl[13429], bl[13430], bl[13431], bl[13432], bl[13433], bl[13434], bl[13435], bl[13436], bl[13437], bl[13438], bl[13439], bl[13440], bl[13441], bl[13442], bl[13443], bl[13444], bl[13445], bl[13446], bl[13447], bl[13448], bl[13449], bl[13450], bl[13451], bl[13452], bl[13453], bl[13454], bl[13455], bl[13456], bl[13457], bl[13458], bl[13459], bl[13460], bl[13461], bl[13462], bl[13463], bl[13464], bl[13465], bl[13466], bl[13467], bl[13468], bl[13469], bl[13470], bl[13471], bl[13472], bl[13473], bl[13474], bl[13475], bl[13476], bl[13477], bl[13478], bl[13479], bl[13480], bl[13481], bl[13482], bl[13483], bl[13484], bl[13485], bl[13486], bl[13487], bl[13488], bl[13489], bl[13490], bl[13491], bl[13492], bl[13493], bl[13494], bl[13495], bl[13496], bl[13497], bl[13498], bl[13499], bl[13500], bl[13501], bl[13502], bl[13503], bl[13504], bl[13505], bl[13506], bl[13507], bl[13508], bl[13509], bl[13510], bl[13511], bl[13512], bl[13513], bl[13514], bl[13515], bl[13516], bl[13517], bl[13518], bl[13519], bl[13520], bl[13521], bl[13522], bl[13523], bl[13524], bl[13525], bl[13526], bl[13527], bl[13528], bl[13529], bl[13530], bl[13531], bl[13532], bl[13533], bl[13534], bl[13535], bl[13536], bl[13537], bl[13538], bl[13539], bl[13540], bl[13541], bl[13542], bl[13543], bl[13544], bl[13545], bl[13546], bl[13547], bl[13548], bl[13549], bl[13550], bl[13551], bl[13552], bl[13553], bl[13554], bl[13555], bl[13556], bl[13557], bl[13558], bl[13559], bl[13560], bl[13561], bl[13562], bl[13563], bl[13564], bl[13565], bl[13566], bl[13567], bl[13568], bl[13569], bl[13570], bl[13571], bl[13572], bl[13573], bl[13574], bl[13575], bl[13576], bl[13577], bl[13578], bl[13579], bl[13580], bl[13581], bl[13582], bl[13583], bl[13584], bl[13585], bl[13586], bl[13587], bl[13588], bl[13589], bl[13590], bl[13591], bl[13592], bl[13593], bl[13594], bl[13595], bl[13596], bl[13597], bl[13598], bl[13599], bl[13600], bl[13601], bl[13602], bl[13603], bl[13604], bl[13605], bl[13606], bl[13607], bl[13608], bl[13609], bl[13610], bl[13611], bl[13612], bl[13613], bl[13614], bl[13615], bl[13616], bl[13617], bl[13618], bl[13619], bl[13620], bl[13621], bl[13622], bl[13623], bl[13624], bl[13625], bl[13626], bl[13627], bl[13628], bl[13629], bl[13630], bl[13631], bl[13632], bl[13633], bl[13634], bl[13635], bl[13636], bl[13637], bl[13638], bl[13639], bl[13640], bl[13641], bl[13642], bl[13643], bl[13644], bl[13645], bl[13646], bl[13647], bl[13648], bl[13649], bl[13650], bl[13651], bl[13652], bl[13653], bl[13654], bl[13655], bl[13656], bl[13657], bl[13658], bl[13659], bl[13660], bl[13661], bl[13662], bl[13663], bl[13664], bl[13665], bl[13666], bl[13667], bl[13668], bl[13669], bl[13670], bl[13671], bl[13672], bl[13673], bl[13674], bl[13675], bl[13676], bl[13677], bl[13678], bl[13679], bl[13680], bl[13681], bl[13682], bl[13683], bl[13684], bl[13685], bl[13686], bl[13687], bl[13688], bl[13689], bl[13690], bl[13691], bl[13692], bl[13693], bl[13694], bl[13695], bl[13696], bl[13697], bl[13698], bl[13699], bl[13700], bl[13701], bl[13702], bl[13703], bl[13704], bl[13705], bl[13706], bl[13707], bl[13708], bl[13709], bl[13710], bl[13711], bl[13712], bl[13713], bl[13714], bl[13715], bl[13716], bl[13717], bl[13718], bl[13719], bl[13720], bl[13721], bl[13722], bl[13723], bl[13724], bl[13725], bl[13726], bl[13727], bl[13728], bl[13729], bl[13730], bl[13731], bl[13732], bl[13733], bl[13734], bl[13735], bl[13736], bl[13737], bl[13738], bl[13739], bl[13740], bl[13741], bl[13742], bl[13743], bl[13744], bl[13745], bl[13746], bl[13747], bl[13748], bl[13749], bl[13750], bl[13751], bl[13752], bl[13753], bl[13754], bl[13755], bl[13756], bl[13757], bl[13758], bl[13759], bl[13760], bl[13761], bl[13762], bl[13763], bl[13764], bl[13765], bl[13766], bl[13767], bl[13768], bl[13769], bl[13770], bl[13771], bl[13772], bl[13773], bl[13774], bl[13775], bl[13776], bl[13777], bl[13778], bl[13779], bl[13780], bl[13781], bl[13782], bl[13783], bl[13784], bl[13785], bl[13786], bl[13787], bl[13788], bl[13789], bl[13790], bl[13791], bl[13792], bl[13793], bl[13794], bl[13795], bl[13796], bl[13797], bl[13798], bl[13799], bl[13800], bl[13801], bl[13802], bl[13803], bl[13804], bl[13805], bl[13806], bl[13807], bl[13808], bl[13809], bl[13810], bl[13811], bl[13812], bl[13813], bl[13814], bl[13815], bl[13816], bl[13817], bl[13818], bl[13819], bl[13820], bl[13821], bl[13822], bl[13823], bl[13824], bl[13825], bl[13826], bl[13827], bl[13828], bl[13829], bl[13830], bl[13831], bl[13832], bl[13833], bl[13834], bl[13835], bl[13836], bl[13837], bl[13838], bl[13839], bl[13840], bl[13841], bl[13842], bl[13843], bl[13844], bl[13845], bl[13846], bl[13847], bl[13848], bl[13849], bl[13850], bl[13851], bl[13852], bl[13853], bl[13854], bl[13855], bl[13856], bl[13857], bl[13858], bl[13859], bl[13860], bl[13861], bl[13862], bl[13863], bl[13864], bl[13865], bl[13866], bl[13867], bl[13868], bl[13869], bl[13870], bl[13871], bl[13872], bl[13873], bl[13874], bl[13875], bl[13876], bl[13877], bl[13878], bl[13879], bl[13880], bl[13881], bl[13882], bl[13883], bl[13884], bl[13885], bl[13886], bl[13887], bl[13888], bl[13889], bl[13890], bl[13891], bl[13892], bl[13893], bl[13894], bl[13895], bl[13896], bl[13897], bl[13898], bl[13899], bl[13900], bl[13901], bl[13902], bl[13903], bl[13904], bl[13905], bl[13906], bl[13907], bl[13908], bl[13909], bl[13910], bl[13911], bl[13912], bl[13913], bl[13914], bl[13915], bl[13916], bl[13917], bl[13918], bl[13919], bl[13920], bl[13921], bl[13922], bl[13923], bl[13924], bl[13925], bl[13926], bl[13927], bl[13928], bl[13929], bl[13930], bl[13931], bl[13932], bl[13933], bl[13934], bl[13935], bl[13936], bl[13937], bl[13938], bl[13939], bl[13940], bl[13941], bl[13942], bl[13943], bl[13944], bl[13945], bl[13946], bl[13947], bl[13948], bl[13949], bl[13950], bl[13951], bl[13952], bl[13953], bl[13954], bl[13955], bl[13956], bl[13957], bl[13958], bl[13959], bl[13960], bl[13961], bl[13962], bl[13963], bl[19068], bl[19069], bl[19070], bl[19071], bl[19072], bl[19073], bl[19074], bl[19075], bl[19076], bl[19077], bl[19078], bl[19079], bl[19080], bl[19081], bl[19082], bl[19083], bl[19084], bl[19085], bl[19086], bl[19087], bl[19088], bl[19089], bl[19090], bl[19091], bl[19092], bl[19093], bl[19094], bl[19095], bl[19096], bl[19097], bl[19098], bl[19099], bl[19100], bl[19101], bl[19102], bl[19103], bl[19104], bl[19105], bl[19106], bl[19107], bl[19108], bl[19109], bl[19110], bl[19111], bl[19112], bl[19113], bl[19114], bl[19115], bl[19116], bl[19117], bl[19118], bl[19119], bl[19120], bl[19121], bl[19122], bl[19123], bl[19124], bl[19125], bl[19126], bl[19127], bl[19128], bl[19129], bl[19130], bl[19131], bl[19132], bl[19133], bl[19134], bl[19135], bl[19136], bl[19137], bl[19138], bl[19139], bl[19140], bl[19141], bl[19142], bl[19143], bl[19144], bl[19145], bl[19146], bl[19147], bl[12864], bl[12865], bl[12866], bl[12867], bl[12868], bl[12869], bl[12870], bl[12871], bl[12872], bl[12873], bl[12874], bl[12875], bl[12876], bl[12877], bl[12878], bl[12879], bl[12880], bl[12881], bl[12882], bl[12883], bl[12884], bl[12885], bl[12886], bl[12887], bl[12888], bl[12889], bl[12890], bl[12891], bl[12892], bl[12893], bl[12894], bl[12895], bl[12896], bl[12897], bl[12898], bl[12899], bl[12900], bl[12901], bl[12902], bl[12903], bl[12904], bl[12905], bl[12906], bl[12907], bl[12908], bl[12909], bl[12910], bl[12911], bl[12912], bl[12913], bl[12914], bl[12915], bl[12916], bl[12917], bl[12918], bl[12919], bl[12920], bl[12921], bl[12922], bl[12923], bl[12924], bl[12925], bl[12926], bl[12927], bl[12928], bl[12929], bl[12930], bl[12931], bl[12932], bl[12933], bl[12934], bl[12935], bl[12936], bl[12937], bl[12938], bl[12939], bl[12940], bl[12941], bl[12942], bl[12943], bl[18988], bl[18989], bl[18990], bl[18991], bl[18992], bl[18993], bl[18994], bl[18995], bl[18996], bl[18997], bl[18998], bl[18999], bl[19000], bl[19001], bl[19002], bl[19003], bl[19004], bl[19005], bl[19006], bl[19007], bl[19008], bl[19009], bl[19010], bl[19011], bl[19012], bl[19013], bl[19014], bl[19015], bl[19016], bl[19017], bl[19018], bl[19019], bl[19020], bl[19021], bl[19022], bl[19023], bl[19024], bl[19025], bl[19026], bl[19027], bl[19028], bl[19029], bl[19030], bl[19031], bl[19032], bl[19033], bl[19034], bl[19035], bl[19036], bl[19037], bl[19038], bl[19039], bl[19040], bl[19041], bl[19042], bl[19043], bl[19044], bl[19045], bl[19046], bl[19047], bl[19048], bl[19049], bl[19050], bl[19051], bl[19052], bl[19053], bl[19054], bl[19055], bl[19056], bl[19057], bl[19058], bl[19059], bl[19060], bl[19061], bl[19062], bl[19063], bl[19064], bl[19065], bl[19066], bl[19067]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    tile tile_4__2_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_2__1__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_2__1__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_2__1__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_3__0__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_3__0__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_3__0__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_2__0__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_2__0__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_2__0__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_2__0__grid_top_r_in[1]),
        .grid_left_in(grid_clb_3__1__grid_left_in),
        .grid_bottom_in(grid_clb_3__1__grid_bottom_in),
        .chanx_left_in(sb_1__1__3_chanx_right_out),
        .chanx_left_out(cbx_1__1__6_chanx_left_out),
        .grid_top_out(grid_clb_3__2__grid_bottom_in),
        .chany_bottom_in(sb_1__0__2_chany_top_out),
        .chany_bottom_out(cby_1__1__8_chany_bottom_out),
        .grid_right_out(grid_clb_4__1__grid_left_in),
        .chany_top_in_0(cby_1__1__9_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__9_chanx_left_out),
        .chany_top_out_0(sb_1__1__6_chany_top_out),
        .chanx_right_out_0(sb_1__1__6_chanx_right_out),
        .grid_top_r_in(sb_3__1__grid_top_r_in),
        .grid_top_l_in(sb_3__1__grid_top_l_in),
        .grid_right_t_in(sb_3__1__grid_right_t_in),
        .grid_right_b_in(sb_3__1__grid_right_b_in),
        .grid_bottom_r_in(sb_3__0__grid_top_r_in),
        .grid_bottom_l_in(sb_3__0__grid_top_l_in),
        .grid_left_t_in(sb_2__1__grid_right_t_in),
        .grid_left_b_in(sb_2__1__grid_right_b_in),
        .bl({bl[4148], bl[4149], bl[4150], bl[4151], bl[4152], bl[4153], bl[4154], bl[4155], bl[4156], bl[4157], bl[4158], bl[4159], bl[4160], bl[4161], bl[4162], bl[4163], bl[4164], bl[4165], bl[4166], bl[4167], bl[4168], bl[4169], bl[4170], bl[4171], bl[4172], bl[4173], bl[4174], bl[4175], bl[4176], bl[4177], bl[4178], bl[4179], bl[4180], bl[4181], bl[4182], bl[4183], bl[4184], bl[4185], bl[4186], bl[4187], bl[4188], bl[4189], bl[4190], bl[4191], bl[4192], bl[4193], bl[4194], bl[4195], bl[4196], bl[4197], bl[4198], bl[4199], bl[4200], bl[4201], bl[4202], bl[4203], bl[4204], bl[4205], bl[4206], bl[4207], bl[4208], bl[4209], bl[4210], bl[4211], bl[4212], bl[4213], bl[4214], bl[4215], bl[4216], bl[4217], bl[4218], bl[4219], bl[4220], bl[4221], bl[4222], bl[4223], bl[4224], bl[4225], bl[4226], bl[4227], bl[4228], bl[4229], bl[4230], bl[4231], bl[4232], bl[4233], bl[4234], bl[4235], bl[4236], bl[4237], bl[4238], bl[4239], bl[4240], bl[4241], bl[4242], bl[4243], bl[4244], bl[4245], bl[4246], bl[4247], bl[4248], bl[4249], bl[4250], bl[4251], bl[4252], bl[4253], bl[4254], bl[4255], bl[4256], bl[4257], bl[4258], bl[4259], bl[4260], bl[4261], bl[4262], bl[4263], bl[4264], bl[4265], bl[4266], bl[4267], bl[4268], bl[4269], bl[4270], bl[4271], bl[4272], bl[4273], bl[4274], bl[4275], bl[4276], bl[4277], bl[4278], bl[4279], bl[4280], bl[4281], bl[4282], bl[4283], bl[4284], bl[4285], bl[4286], bl[4287], bl[4288], bl[4289], bl[4290], bl[4291], bl[4292], bl[4293], bl[4294], bl[4295], bl[4296], bl[4297], bl[4298], bl[4299], bl[4300], bl[4301], bl[4302], bl[4303], bl[4304], bl[4305], bl[4306], bl[4307], bl[4308], bl[4309], bl[4310], bl[4311], bl[4312], bl[4313], bl[4314], bl[4315], bl[4316], bl[4317], bl[4318], bl[4319], bl[4320], bl[4321], bl[4322], bl[4323], bl[4324], bl[4325], bl[4326], bl[4327], bl[4328], bl[4329], bl[4330], bl[4331], bl[4332], bl[4333], bl[4334], bl[4335], bl[4336], bl[4337], bl[4338], bl[4339], bl[4340], bl[4341], bl[4342], bl[4343], bl[4344], bl[4345], bl[4346], bl[4347], bl[4348], bl[4349], bl[4350], bl[4351], bl[4352], bl[4353], bl[4354], bl[4355], bl[4356], bl[4357], bl[4358], bl[4359], bl[4360], bl[4361], bl[4362], bl[4363], bl[4364], bl[4365], bl[4366], bl[4367], bl[4368], bl[4369], bl[4370], bl[4371], bl[4372], bl[4373], bl[4374], bl[4375], bl[4376], bl[4377], bl[4378], bl[4379], bl[4380], bl[4381], bl[4382], bl[4383], bl[4384], bl[4385], bl[4386], bl[4387], bl[4388], bl[4389], bl[4390], bl[4391], bl[4392], bl[4393], bl[4394], bl[4395], bl[4396], bl[4397], bl[4398], bl[4399], bl[4400], bl[4401], bl[4402], bl[4403], bl[4404], bl[4405], bl[4406], bl[4407], bl[4408], bl[4409], bl[4410], bl[4411], bl[4412], bl[4413], bl[4414], bl[4415], bl[4416], bl[4417], bl[4418], bl[4419], bl[4420], bl[4421], bl[4422], bl[4423], bl[4424], bl[4425], bl[4426], bl[4427], bl[4428], bl[4429], bl[4430], bl[4431], bl[4432], bl[4433], bl[4434], bl[4435], bl[4436], bl[4437], bl[4438], bl[4439], bl[4440], bl[4441], bl[4442], bl[4443], bl[4444], bl[4445], bl[4446], bl[4447], bl[4448], bl[4449], bl[4450], bl[4451], bl[4452], bl[4453], bl[4454], bl[4455], bl[4456], bl[4457], bl[4458], bl[4459], bl[4460], bl[4461], bl[4462], bl[4463], bl[4464], bl[4465], bl[4466], bl[4467], bl[4468], bl[4469], bl[4470], bl[4471], bl[4472], bl[4473], bl[4474], bl[4475], bl[4476], bl[4477], bl[4478], bl[4479], bl[4480], bl[4481], bl[4482], bl[4483], bl[4484], bl[4485], bl[4486], bl[4487], bl[4488], bl[4489], bl[4490], bl[4491], bl[4492], bl[4493], bl[4494], bl[4495], bl[4496], bl[4497], bl[4498], bl[4499], bl[4500], bl[4501], bl[4502], bl[4503], bl[4504], bl[4505], bl[4506], bl[4507], bl[4508], bl[4509], bl[4510], bl[4511], bl[4512], bl[4513], bl[4514], bl[4515], bl[4516], bl[4517], bl[4518], bl[4519], bl[4520], bl[4521], bl[4522], bl[4523], bl[4524], bl[4525], bl[4526], bl[4527], bl[4528], bl[4529], bl[4530], bl[4531], bl[4532], bl[4533], bl[4534], bl[4535], bl[4536], bl[4537], bl[4538], bl[4539], bl[4540], bl[4541], bl[4542], bl[4543], bl[4544], bl[4545], bl[4546], bl[4547], bl[4548], bl[4549], bl[4550], bl[4551], bl[4552], bl[4553], bl[4554], bl[4555], bl[4556], bl[4557], bl[4558], bl[4559], bl[4560], bl[4561], bl[4562], bl[4563], bl[4564], bl[4565], bl[4566], bl[4567], bl[4568], bl[4569], bl[4570], bl[4571], bl[4572], bl[4573], bl[4574], bl[4575], bl[4576], bl[4577], bl[4578], bl[4579], bl[4580], bl[4581], bl[4582], bl[4583], bl[4584], bl[4585], bl[4586], bl[4587], bl[4588], bl[4589], bl[4590], bl[4591], bl[4592], bl[4593], bl[4594], bl[4595], bl[4596], bl[4597], bl[4598], bl[4599], bl[4600], bl[4601], bl[4602], bl[4603], bl[4604], bl[4605], bl[4606], bl[4607], bl[4608], bl[4609], bl[4610], bl[4611], bl[4612], bl[4613], bl[4614], bl[4615], bl[4616], bl[4617], bl[4618], bl[4619], bl[4620], bl[4621], bl[4622], bl[4623], bl[4624], bl[4625], bl[4626], bl[4627], bl[4628], bl[4629], bl[4630], bl[4631], bl[4632], bl[4633], bl[4634], bl[4635], bl[4636], bl[4637], bl[4638], bl[4639], bl[4640], bl[4641], bl[4642], bl[4643], bl[4644], bl[4645], bl[4646], bl[4647], bl[4648], bl[4649], bl[4650], bl[4651], bl[4652], bl[4653], bl[4654], bl[4655], bl[4656], bl[4657], bl[4658], bl[4659], bl[4660], bl[4661], bl[4662], bl[4663], bl[4664], bl[4665], bl[4666], bl[4667], bl[4668], bl[4669], bl[4670], bl[4671], bl[4672], bl[4673], bl[4674], bl[4675], bl[4676], bl[4677], bl[4678], bl[4679], bl[4680], bl[4681], bl[4682], bl[4683], bl[4684], bl[4685], bl[4686], bl[4687], bl[4688], bl[4689], bl[4690], bl[4691], bl[4692], bl[4693], bl[4694], bl[4695], bl[4696], bl[4697], bl[4698], bl[4699], bl[4700], bl[4701], bl[4702], bl[4703], bl[4704], bl[4705], bl[4706], bl[4707], bl[4708], bl[4709], bl[4710], bl[4711], bl[4712], bl[4713], bl[4714], bl[4715], bl[4716], bl[4717], bl[4718], bl[4719], bl[4720], bl[4721], bl[4722], bl[4723], bl[4724], bl[4725], bl[4726], bl[4727], bl[4728], bl[4729], bl[4730], bl[4731], bl[4732], bl[4733], bl[4734], bl[4735], bl[4736], bl[4737], bl[4738], bl[4739], bl[4740], bl[4741], bl[4742], bl[4743], bl[4744], bl[4745], bl[4746], bl[4747], bl[4748], bl[4749], bl[4750], bl[4751], bl[4752], bl[4753], bl[4754], bl[4755], bl[4756], bl[4757], bl[4758], bl[4759], bl[4760], bl[4761], bl[4762], bl[4763], bl[4764], bl[4765], bl[4766], bl[4767], bl[4768], bl[4769], bl[4770], bl[4771], bl[4772], bl[4773], bl[4774], bl[4775], bl[4776], bl[4777], bl[4778], bl[4779], bl[4780], bl[4781], bl[4782], bl[4783], bl[4784], bl[4785], bl[4786], bl[4787], bl[4788], bl[4789], bl[4790], bl[4791], bl[4792], bl[4793], bl[4794], bl[4795], bl[4796], bl[4797], bl[4798], bl[4799], bl[4800], bl[4801], bl[4802], bl[4803], bl[4804], bl[4805], bl[4806], bl[4807], bl[4808], bl[4809], bl[4810], bl[4811], bl[4812], bl[4813], bl[4814], bl[4815], bl[4816], bl[4817], bl[4818], bl[4819], bl[4820], bl[4821], bl[4822], bl[4823], bl[4824], bl[4825], bl[4826], bl[4827], bl[4828], bl[4829], bl[4830], bl[4831], bl[4832], bl[4833], bl[4834], bl[4835], bl[4836], bl[4837], bl[4838], bl[4839], bl[4840], bl[4841], bl[4842], bl[4843], bl[4844], bl[4845], bl[4846], bl[4847], bl[4848], bl[4849], bl[4850], bl[4851], bl[4852], bl[4853], bl[4854], bl[4855], bl[4856], bl[4857], bl[4858], bl[4859], bl[4860], bl[4861], bl[4862], bl[4863], bl[4864], bl[4865], bl[4866], bl[4867], bl[4868], bl[4869], bl[4870], bl[4871], bl[4872], bl[4873], bl[4874], bl[4875], bl[4876], bl[4877], bl[4878], bl[4879], bl[4880], bl[4881], bl[4882], bl[4883], bl[4884], bl[4885], bl[4886], bl[4887], bl[4888], bl[4889], bl[4890], bl[4891], bl[4892], bl[4893], bl[4894], bl[4895], bl[4896], bl[4897], bl[4898], bl[4899], bl[4900], bl[4901], bl[4902], bl[4903], bl[4904], bl[4905], bl[4906], bl[4907], bl[4908], bl[4909], bl[4910], bl[4911], bl[4912], bl[4913], bl[4914], bl[4915], bl[4916], bl[4917], bl[4918], bl[4919], bl[4920], bl[4921], bl[4922], bl[4923], bl[4924], bl[4925], bl[4926], bl[4927], bl[4928], bl[4929], bl[4930], bl[4931], bl[4932], bl[4933], bl[4934], bl[4935], bl[4936], bl[4937], bl[4938], bl[4939], bl[4940], bl[4941], bl[4942], bl[4943], bl[4944], bl[4945], bl[4946], bl[4947], bl[4948], bl[4949], bl[4950], bl[4951], bl[4952], bl[4953], bl[4954], bl[4955], bl[4956], bl[4957], bl[4958], bl[4959], bl[4960], bl[4961], bl[4962], bl[4963], bl[4964], bl[4965], bl[4966], bl[4967], bl[4968], bl[4969], bl[4970], bl[4971], bl[4972], bl[4973], bl[4974], bl[4975], bl[4976], bl[4977], bl[4978], bl[4979], bl[4980], bl[4981], bl[4982], bl[4983], bl[4984], bl[4985], bl[4986], bl[4987], bl[4988], bl[4989], bl[4990], bl[4991], bl[4992], bl[4993], bl[4994], bl[4995], bl[4996], bl[4997], bl[4998], bl[4999], bl[5000], bl[5001], bl[5002], bl[5003], bl[5004], bl[5005], bl[5006], bl[5007], bl[5008], bl[5009], bl[5010], bl[5011], bl[5012], bl[5013], bl[5014], bl[5015], bl[5016], bl[5017], bl[5018], bl[5019], bl[5020], bl[5021], bl[5022], bl[5023], bl[5024], bl[5025], bl[5026], bl[5027], bl[5028], bl[5029], bl[5030], bl[5031], bl[5032], bl[5033], bl[5034], bl[5035], bl[5036], bl[5037], bl[5038], bl[5039], bl[5040], bl[5041], bl[5042], bl[5043], bl[5044], bl[5045], bl[5046], bl[5047], bl[5048], bl[5049], bl[5050], bl[5051], bl[5052], bl[5053], bl[5054], bl[5055], bl[5056], bl[5057], bl[5058], bl[5059], bl[5060], bl[5061], bl[5062], bl[5063], bl[5064], bl[5065], bl[5066], bl[5067], bl[5068], bl[5069], bl[5070], bl[5071], bl[5072], bl[5073], bl[5074], bl[5075], bl[5076], bl[5077], bl[5078], bl[5079], bl[5080], bl[5081], bl[5082], bl[5083], bl[5084], bl[5085], bl[5086], bl[5087], bl[5088], bl[5089], bl[5090], bl[5091], bl[5092], bl[5093], bl[5094], bl[5095], bl[5096], bl[5097], bl[5098], bl[5099], bl[5100], bl[5101], bl[5102], bl[5103], bl[5104], bl[5105], bl[5106], bl[5107], bl[5108], bl[5109], bl[5110], bl[5111], bl[5112], bl[5113], bl[5114], bl[5115], bl[5116], bl[5117], bl[5118], bl[5119], bl[5120], bl[5121], bl[5122], bl[5123], bl[5124], bl[5125], bl[5126], bl[5127], bl[5128], bl[5129], bl[5130], bl[5131], bl[5132], bl[5133], bl[5134], bl[5135], bl[5136], bl[5137], bl[5138], bl[5139], bl[5140], bl[5141], bl[5142], bl[5143], bl[5144], bl[5145], bl[5146], bl[5147], bl[5148], bl[5149], bl[5150], bl[5151], bl[5152], bl[5153], bl[5154], bl[5155], bl[5156], bl[5157], bl[5158], bl[5159], bl[5160], bl[5161], bl[5162], bl[5163], bl[5164], bl[5165], bl[5166], bl[5167], bl[7744], bl[7745], bl[7746], bl[7747], bl[7748], bl[7749], bl[7750], bl[7751], bl[7752], bl[7753], bl[7754], bl[7755], bl[7756], bl[7757], bl[7758], bl[7759], bl[7760], bl[7761], bl[7762], bl[7763], bl[7764], bl[7765], bl[7766], bl[7767], bl[7768], bl[7769], bl[7770], bl[7771], bl[7772], bl[7773], bl[7774], bl[7775], bl[7776], bl[7777], bl[7778], bl[7779], bl[7780], bl[7781], bl[7782], bl[7783], bl[7784], bl[7785], bl[7786], bl[7787], bl[7788], bl[7789], bl[7790], bl[7791], bl[7792], bl[7793], bl[7794], bl[7795], bl[7796], bl[7797], bl[7798], bl[7799], bl[7800], bl[7801], bl[7802], bl[7803], bl[7804], bl[7805], bl[7806], bl[7807], bl[7808], bl[7809], bl[7810], bl[7811], bl[7812], bl[7813], bl[7814], bl[7815], bl[7816], bl[7817], bl[7818], bl[7819], bl[7820], bl[7821], bl[7822], bl[7823], bl[4068], bl[4069], bl[4070], bl[4071], bl[4072], bl[4073], bl[4074], bl[4075], bl[4076], bl[4077], bl[4078], bl[4079], bl[4080], bl[4081], bl[4082], bl[4083], bl[4084], bl[4085], bl[4086], bl[4087], bl[4088], bl[4089], bl[4090], bl[4091], bl[4092], bl[4093], bl[4094], bl[4095], bl[4096], bl[4097], bl[4098], bl[4099], bl[4100], bl[4101], bl[4102], bl[4103], bl[4104], bl[4105], bl[4106], bl[4107], bl[4108], bl[4109], bl[4110], bl[4111], bl[4112], bl[4113], bl[4114], bl[4115], bl[4116], bl[4117], bl[4118], bl[4119], bl[4120], bl[4121], bl[4122], bl[4123], bl[4124], bl[4125], bl[4126], bl[4127], bl[4128], bl[4129], bl[4130], bl[4131], bl[4132], bl[4133], bl[4134], bl[4135], bl[4136], bl[4137], bl[4138], bl[4139], bl[4140], bl[4141], bl[4142], bl[4143], bl[4144], bl[4145], bl[4146], bl[4147], bl[7664], bl[7665], bl[7666], bl[7667], bl[7668], bl[7669], bl[7670], bl[7671], bl[7672], bl[7673], bl[7674], bl[7675], bl[7676], bl[7677], bl[7678], bl[7679], bl[7680], bl[7681], bl[7682], bl[7683], bl[7684], bl[7685], bl[7686], bl[7687], bl[7688], bl[7689], bl[7690], bl[7691], bl[7692], bl[7693], bl[7694], bl[7695], bl[7696], bl[7697], bl[7698], bl[7699], bl[7700], bl[7701], bl[7702], bl[7703], bl[7704], bl[7705], bl[7706], bl[7707], bl[7708], bl[7709], bl[7710], bl[7711], bl[7712], bl[7713], bl[7714], bl[7715], bl[7716], bl[7717], bl[7718], bl[7719], bl[7720], bl[7721], bl[7722], bl[7723], bl[7724], bl[7725], bl[7726], bl[7727], bl[7728], bl[7729], bl[7730], bl[7731], bl[7732], bl[7733], bl[7734], bl[7735], bl[7736], bl[7737], bl[7738], bl[7739], bl[7740], bl[7741], bl[7742], bl[7743]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    tile tile_4__3_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_2__2__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_2__2__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_2__2__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_3__1__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_3__1__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_3__1__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_2__1__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_2__1__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_2__1__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_2__1__grid_top_r_in[1]),
        .grid_left_in(grid_clb_3__2__grid_left_in),
        .grid_bottom_in(grid_clb_3__2__grid_bottom_in),
        .chanx_left_in(sb_1__1__4_chanx_right_out),
        .chanx_left_out(cbx_1__1__7_chanx_left_out),
        .grid_top_out(grid_clb_3__3__grid_bottom_in),
        .chany_bottom_in(sb_1__1__6_chany_top_out),
        .chany_bottom_out(cby_1__1__9_chany_bottom_out),
        .grid_right_out(grid_clb_4__2__grid_left_in),
        .chany_top_in_0(cby_1__1__10_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__10_chanx_left_out),
        .chany_top_out_0(sb_1__1__7_chany_top_out),
        .chanx_right_out_0(sb_1__1__7_chanx_right_out),
        .grid_top_r_in(sb_3__2__grid_top_r_in),
        .grid_top_l_in(sb_3__2__grid_top_l_in),
        .grid_right_t_in(sb_3__2__grid_right_t_in),
        .grid_right_b_in(sb_3__2__grid_right_b_in),
        .grid_bottom_r_in(sb_3__1__grid_top_r_in),
        .grid_bottom_l_in(sb_3__1__grid_top_l_in),
        .grid_left_t_in(sb_2__2__grid_right_t_in),
        .grid_left_b_in(sb_2__2__grid_right_b_in),
        .bl({bl[7904], bl[7905], bl[7906], bl[7907], bl[7908], bl[7909], bl[7910], bl[7911], bl[7912], bl[7913], bl[7914], bl[7915], bl[7916], bl[7917], bl[7918], bl[7919], bl[7920], bl[7921], bl[7922], bl[7923], bl[7924], bl[7925], bl[7926], bl[7927], bl[7928], bl[7929], bl[7930], bl[7931], bl[7932], bl[7933], bl[7934], bl[7935], bl[7936], bl[7937], bl[7938], bl[7939], bl[7940], bl[7941], bl[7942], bl[7943], bl[7944], bl[7945], bl[7946], bl[7947], bl[7948], bl[7949], bl[7950], bl[7951], bl[7952], bl[7953], bl[7954], bl[7955], bl[7956], bl[7957], bl[7958], bl[7959], bl[7960], bl[7961], bl[7962], bl[7963], bl[7964], bl[7965], bl[7966], bl[7967], bl[7968], bl[7969], bl[7970], bl[7971], bl[7972], bl[7973], bl[7974], bl[7975], bl[7976], bl[7977], bl[7978], bl[7979], bl[7980], bl[7981], bl[7982], bl[7983], bl[7984], bl[7985], bl[7986], bl[7987], bl[7988], bl[7989], bl[7990], bl[7991], bl[7992], bl[7993], bl[7994], bl[7995], bl[7996], bl[7997], bl[7998], bl[7999], bl[8000], bl[8001], bl[8002], bl[8003], bl[8004], bl[8005], bl[8006], bl[8007], bl[8008], bl[8009], bl[8010], bl[8011], bl[8012], bl[8013], bl[8014], bl[8015], bl[8016], bl[8017], bl[8018], bl[8019], bl[8020], bl[8021], bl[8022], bl[8023], bl[8024], bl[8025], bl[8026], bl[8027], bl[8028], bl[8029], bl[8030], bl[8031], bl[8032], bl[8033], bl[8034], bl[8035], bl[8036], bl[8037], bl[8038], bl[8039], bl[8040], bl[8041], bl[8042], bl[8043], bl[8044], bl[8045], bl[8046], bl[8047], bl[8048], bl[8049], bl[8050], bl[8051], bl[8052], bl[8053], bl[8054], bl[8055], bl[8056], bl[8057], bl[8058], bl[8059], bl[8060], bl[8061], bl[8062], bl[8063], bl[8064], bl[8065], bl[8066], bl[8067], bl[8068], bl[8069], bl[8070], bl[8071], bl[8072], bl[8073], bl[8074], bl[8075], bl[8076], bl[8077], bl[8078], bl[8079], bl[8080], bl[8081], bl[8082], bl[8083], bl[8084], bl[8085], bl[8086], bl[8087], bl[8088], bl[8089], bl[8090], bl[8091], bl[8092], bl[8093], bl[8094], bl[8095], bl[8096], bl[8097], bl[8098], bl[8099], bl[8100], bl[8101], bl[8102], bl[8103], bl[8104], bl[8105], bl[8106], bl[8107], bl[8108], bl[8109], bl[8110], bl[8111], bl[8112], bl[8113], bl[8114], bl[8115], bl[8116], bl[8117], bl[8118], bl[8119], bl[8120], bl[8121], bl[8122], bl[8123], bl[8124], bl[8125], bl[8126], bl[8127], bl[8128], bl[8129], bl[8130], bl[8131], bl[8132], bl[8133], bl[8134], bl[8135], bl[8136], bl[8137], bl[8138], bl[8139], bl[8140], bl[8141], bl[8142], bl[8143], bl[8144], bl[8145], bl[8146], bl[8147], bl[8148], bl[8149], bl[8150], bl[8151], bl[8152], bl[8153], bl[8154], bl[8155], bl[8156], bl[8157], bl[8158], bl[8159], bl[8160], bl[8161], bl[8162], bl[8163], bl[8164], bl[8165], bl[8166], bl[8167], bl[8168], bl[8169], bl[8170], bl[8171], bl[8172], bl[8173], bl[8174], bl[8175], bl[8176], bl[8177], bl[8178], bl[8179], bl[8180], bl[8181], bl[8182], bl[8183], bl[8184], bl[8185], bl[8186], bl[8187], bl[8188], bl[8189], bl[8190], bl[8191], bl[8192], bl[8193], bl[8194], bl[8195], bl[8196], bl[8197], bl[8198], bl[8199], bl[8200], bl[8201], bl[8202], bl[8203], bl[8204], bl[8205], bl[8206], bl[8207], bl[8208], bl[8209], bl[8210], bl[8211], bl[8212], bl[8213], bl[8214], bl[8215], bl[8216], bl[8217], bl[8218], bl[8219], bl[8220], bl[8221], bl[8222], bl[8223], bl[8224], bl[8225], bl[8226], bl[8227], bl[8228], bl[8229], bl[8230], bl[8231], bl[8232], bl[8233], bl[8234], bl[8235], bl[8236], bl[8237], bl[8238], bl[8239], bl[8240], bl[8241], bl[8242], bl[8243], bl[8244], bl[8245], bl[8246], bl[8247], bl[8248], bl[8249], bl[8250], bl[8251], bl[8252], bl[8253], bl[8254], bl[8255], bl[8256], bl[8257], bl[8258], bl[8259], bl[8260], bl[8261], bl[8262], bl[8263], bl[8264], bl[8265], bl[8266], bl[8267], bl[8268], bl[8269], bl[8270], bl[8271], bl[8272], bl[8273], bl[8274], bl[8275], bl[8276], bl[8277], bl[8278], bl[8279], bl[8280], bl[8281], bl[8282], bl[8283], bl[8284], bl[8285], bl[8286], bl[8287], bl[8288], bl[8289], bl[8290], bl[8291], bl[8292], bl[8293], bl[8294], bl[8295], bl[8296], bl[8297], bl[8298], bl[8299], bl[8300], bl[8301], bl[8302], bl[8303], bl[8304], bl[8305], bl[8306], bl[8307], bl[8308], bl[8309], bl[8310], bl[8311], bl[8312], bl[8313], bl[8314], bl[8315], bl[8316], bl[8317], bl[8318], bl[8319], bl[8320], bl[8321], bl[8322], bl[8323], bl[8324], bl[8325], bl[8326], bl[8327], bl[8328], bl[8329], bl[8330], bl[8331], bl[8332], bl[8333], bl[8334], bl[8335], bl[8336], bl[8337], bl[8338], bl[8339], bl[8340], bl[8341], bl[8342], bl[8343], bl[8344], bl[8345], bl[8346], bl[8347], bl[8348], bl[8349], bl[8350], bl[8351], bl[8352], bl[8353], bl[8354], bl[8355], bl[8356], bl[8357], bl[8358], bl[8359], bl[8360], bl[8361], bl[8362], bl[8363], bl[8364], bl[8365], bl[8366], bl[8367], bl[8368], bl[8369], bl[8370], bl[8371], bl[8372], bl[8373], bl[8374], bl[8375], bl[8376], bl[8377], bl[8378], bl[8379], bl[8380], bl[8381], bl[8382], bl[8383], bl[8384], bl[8385], bl[8386], bl[8387], bl[8388], bl[8389], bl[8390], bl[8391], bl[8392], bl[8393], bl[8394], bl[8395], bl[8396], bl[8397], bl[8398], bl[8399], bl[8400], bl[8401], bl[8402], bl[8403], bl[8404], bl[8405], bl[8406], bl[8407], bl[8408], bl[8409], bl[8410], bl[8411], bl[8412], bl[8413], bl[8414], bl[8415], bl[8416], bl[8417], bl[8418], bl[8419], bl[8420], bl[8421], bl[8422], bl[8423], bl[8424], bl[8425], bl[8426], bl[8427], bl[8428], bl[8429], bl[8430], bl[8431], bl[8432], bl[8433], bl[8434], bl[8435], bl[8436], bl[8437], bl[8438], bl[8439], bl[8440], bl[8441], bl[8442], bl[8443], bl[8444], bl[8445], bl[8446], bl[8447], bl[8448], bl[8449], bl[8450], bl[8451], bl[8452], bl[8453], bl[8454], bl[8455], bl[8456], bl[8457], bl[8458], bl[8459], bl[8460], bl[8461], bl[8462], bl[8463], bl[8464], bl[8465], bl[8466], bl[8467], bl[8468], bl[8469], bl[8470], bl[8471], bl[8472], bl[8473], bl[8474], bl[8475], bl[8476], bl[8477], bl[8478], bl[8479], bl[8480], bl[8481], bl[8482], bl[8483], bl[8484], bl[8485], bl[8486], bl[8487], bl[8488], bl[8489], bl[8490], bl[8491], bl[8492], bl[8493], bl[8494], bl[8495], bl[8496], bl[8497], bl[8498], bl[8499], bl[8500], bl[8501], bl[8502], bl[8503], bl[8504], bl[8505], bl[8506], bl[8507], bl[8508], bl[8509], bl[8510], bl[8511], bl[8512], bl[8513], bl[8514], bl[8515], bl[8516], bl[8517], bl[8518], bl[8519], bl[8520], bl[8521], bl[8522], bl[8523], bl[8524], bl[8525], bl[8526], bl[8527], bl[8528], bl[8529], bl[8530], bl[8531], bl[8532], bl[8533], bl[8534], bl[8535], bl[8536], bl[8537], bl[8538], bl[8539], bl[8540], bl[8541], bl[8542], bl[8543], bl[8544], bl[8545], bl[8546], bl[8547], bl[8548], bl[8549], bl[8550], bl[8551], bl[8552], bl[8553], bl[8554], bl[8555], bl[8556], bl[8557], bl[8558], bl[8559], bl[8560], bl[8561], bl[8562], bl[8563], bl[8564], bl[8565], bl[8566], bl[8567], bl[8568], bl[8569], bl[8570], bl[8571], bl[8572], bl[8573], bl[8574], bl[8575], bl[8576], bl[8577], bl[8578], bl[8579], bl[8580], bl[8581], bl[8582], bl[8583], bl[8584], bl[8585], bl[8586], bl[8587], bl[8588], bl[8589], bl[8590], bl[8591], bl[8592], bl[8593], bl[8594], bl[8595], bl[8596], bl[8597], bl[8598], bl[8599], bl[8600], bl[8601], bl[8602], bl[8603], bl[8604], bl[8605], bl[8606], bl[8607], bl[8608], bl[8609], bl[8610], bl[8611], bl[8612], bl[8613], bl[8614], bl[8615], bl[8616], bl[8617], bl[8618], bl[8619], bl[8620], bl[8621], bl[8622], bl[8623], bl[8624], bl[8625], bl[8626], bl[8627], bl[8628], bl[8629], bl[8630], bl[8631], bl[8632], bl[8633], bl[8634], bl[8635], bl[8636], bl[8637], bl[8638], bl[8639], bl[8640], bl[8641], bl[8642], bl[8643], bl[8644], bl[8645], bl[8646], bl[8647], bl[8648], bl[8649], bl[8650], bl[8651], bl[8652], bl[8653], bl[8654], bl[8655], bl[8656], bl[8657], bl[8658], bl[8659], bl[8660], bl[8661], bl[8662], bl[8663], bl[8664], bl[8665], bl[8666], bl[8667], bl[8668], bl[8669], bl[8670], bl[8671], bl[8672], bl[8673], bl[8674], bl[8675], bl[8676], bl[8677], bl[8678], bl[8679], bl[8680], bl[8681], bl[8682], bl[8683], bl[8684], bl[8685], bl[8686], bl[8687], bl[8688], bl[8689], bl[8690], bl[8691], bl[8692], bl[8693], bl[8694], bl[8695], bl[8696], bl[8697], bl[8698], bl[8699], bl[8700], bl[8701], bl[8702], bl[8703], bl[8704], bl[8705], bl[8706], bl[8707], bl[8708], bl[8709], bl[8710], bl[8711], bl[8712], bl[8713], bl[8714], bl[8715], bl[8716], bl[8717], bl[8718], bl[8719], bl[8720], bl[8721], bl[8722], bl[8723], bl[8724], bl[8725], bl[8726], bl[8727], bl[8728], bl[8729], bl[8730], bl[8731], bl[8732], bl[8733], bl[8734], bl[8735], bl[8736], bl[8737], bl[8738], bl[8739], bl[8740], bl[8741], bl[8742], bl[8743], bl[8744], bl[8745], bl[8746], bl[8747], bl[8748], bl[8749], bl[8750], bl[8751], bl[8752], bl[8753], bl[8754], bl[8755], bl[8756], bl[8757], bl[8758], bl[8759], bl[8760], bl[8761], bl[8762], bl[8763], bl[8764], bl[8765], bl[8766], bl[8767], bl[8768], bl[8769], bl[8770], bl[8771], bl[8772], bl[8773], bl[8774], bl[8775], bl[8776], bl[8777], bl[8778], bl[8779], bl[8780], bl[8781], bl[8782], bl[8783], bl[8784], bl[8785], bl[8786], bl[8787], bl[8788], bl[8789], bl[8790], bl[8791], bl[8792], bl[8793], bl[8794], bl[8795], bl[8796], bl[8797], bl[8798], bl[8799], bl[8800], bl[8801], bl[8802], bl[8803], bl[8804], bl[8805], bl[8806], bl[8807], bl[8808], bl[8809], bl[8810], bl[8811], bl[8812], bl[8813], bl[8814], bl[8815], bl[8816], bl[8817], bl[8818], bl[8819], bl[8820], bl[8821], bl[8822], bl[8823], bl[8824], bl[8825], bl[8826], bl[8827], bl[8828], bl[8829], bl[8830], bl[8831], bl[8832], bl[8833], bl[8834], bl[8835], bl[8836], bl[8837], bl[8838], bl[8839], bl[8840], bl[8841], bl[8842], bl[8843], bl[8844], bl[8845], bl[8846], bl[8847], bl[8848], bl[8849], bl[8850], bl[8851], bl[8852], bl[8853], bl[8854], bl[8855], bl[8856], bl[8857], bl[8858], bl[8859], bl[8860], bl[8861], bl[8862], bl[8863], bl[8864], bl[8865], bl[8866], bl[8867], bl[8868], bl[8869], bl[8870], bl[8871], bl[8872], bl[8873], bl[8874], bl[8875], bl[8876], bl[8877], bl[8878], bl[8879], bl[8880], bl[8881], bl[8882], bl[8883], bl[8884], bl[8885], bl[8886], bl[8887], bl[8888], bl[8889], bl[8890], bl[8891], bl[8892], bl[8893], bl[8894], bl[8895], bl[8896], bl[8897], bl[8898], bl[8899], bl[8900], bl[8901], bl[8902], bl[8903], bl[8904], bl[8905], bl[8906], bl[8907], bl[8908], bl[8909], bl[8910], bl[8911], bl[8912], bl[8913], bl[8914], bl[8915], bl[8916], bl[8917], bl[8918], bl[8919], bl[8920], bl[8921], bl[8922], bl[8923], bl[14044], bl[14045], bl[14046], bl[14047], bl[14048], bl[14049], bl[14050], bl[14051], bl[14052], bl[14053], bl[14054], bl[14055], bl[14056], bl[14057], bl[14058], bl[14059], bl[14060], bl[14061], bl[14062], bl[14063], bl[14064], bl[14065], bl[14066], bl[14067], bl[14068], bl[14069], bl[14070], bl[14071], bl[14072], bl[14073], bl[14074], bl[14075], bl[14076], bl[14077], bl[14078], bl[14079], bl[14080], bl[14081], bl[14082], bl[14083], bl[14084], bl[14085], bl[14086], bl[14087], bl[14088], bl[14089], bl[14090], bl[14091], bl[14092], bl[14093], bl[14094], bl[14095], bl[14096], bl[14097], bl[14098], bl[14099], bl[14100], bl[14101], bl[14102], bl[14103], bl[14104], bl[14105], bl[14106], bl[14107], bl[14108], bl[14109], bl[14110], bl[14111], bl[14112], bl[14113], bl[14114], bl[14115], bl[14116], bl[14117], bl[14118], bl[14119], bl[14120], bl[14121], bl[14122], bl[14123], bl[7824], bl[7825], bl[7826], bl[7827], bl[7828], bl[7829], bl[7830], bl[7831], bl[7832], bl[7833], bl[7834], bl[7835], bl[7836], bl[7837], bl[7838], bl[7839], bl[7840], bl[7841], bl[7842], bl[7843], bl[7844], bl[7845], bl[7846], bl[7847], bl[7848], bl[7849], bl[7850], bl[7851], bl[7852], bl[7853], bl[7854], bl[7855], bl[7856], bl[7857], bl[7858], bl[7859], bl[7860], bl[7861], bl[7862], bl[7863], bl[7864], bl[7865], bl[7866], bl[7867], bl[7868], bl[7869], bl[7870], bl[7871], bl[7872], bl[7873], bl[7874], bl[7875], bl[7876], bl[7877], bl[7878], bl[7879], bl[7880], bl[7881], bl[7882], bl[7883], bl[7884], bl[7885], bl[7886], bl[7887], bl[7888], bl[7889], bl[7890], bl[7891], bl[7892], bl[7893], bl[7894], bl[7895], bl[7896], bl[7897], bl[7898], bl[7899], bl[7900], bl[7901], bl[7902], bl[7903], bl[13964], bl[13965], bl[13966], bl[13967], bl[13968], bl[13969], bl[13970], bl[13971], bl[13972], bl[13973], bl[13974], bl[13975], bl[13976], bl[13977], bl[13978], bl[13979], bl[13980], bl[13981], bl[13982], bl[13983], bl[13984], bl[13985], bl[13986], bl[13987], bl[13988], bl[13989], bl[13990], bl[13991], bl[13992], bl[13993], bl[13994], bl[13995], bl[13996], bl[13997], bl[13998], bl[13999], bl[14000], bl[14001], bl[14002], bl[14003], bl[14004], bl[14005], bl[14006], bl[14007], bl[14008], bl[14009], bl[14010], bl[14011], bl[14012], bl[14013], bl[14014], bl[14015], bl[14016], bl[14017], bl[14018], bl[14019], bl[14020], bl[14021], bl[14022], bl[14023], bl[14024], bl[14025], bl[14026], bl[14027], bl[14028], bl[14029], bl[14030], bl[14031], bl[14032], bl[14033], bl[14034], bl[14035], bl[14036], bl[14037], bl[14038], bl[14039], bl[14040], bl[14041], bl[14042], bl[14043]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    tile tile_4__4_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_2__3__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_2__3__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_2__3__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_3__2__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_3__2__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_3__2__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_2__2__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_2__2__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_2__2__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_2__2__grid_top_r_in[1]),
        .grid_left_in(grid_clb_3__3__grid_left_in),
        .grid_bottom_in(grid_clb_3__3__grid_bottom_in),
        .chanx_left_in(sb_1__1__5_chanx_right_out),
        .chanx_left_out(cbx_1__1__8_chanx_left_out),
        .grid_top_out(grid_clb_3__4__grid_bottom_in),
        .chany_bottom_in(sb_1__1__7_chany_top_out),
        .chany_bottom_out(cby_1__1__10_chany_bottom_out),
        .grid_right_out(grid_clb_4__3__grid_left_in),
        .chany_top_in_0(cby_1__1__11_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__11_chanx_left_out),
        .chany_top_out_0(sb_1__1__8_chany_top_out),
        .chanx_right_out_0(sb_1__1__8_chanx_right_out),
        .grid_top_r_in(sb_3__3__grid_top_r_in),
        .grid_top_l_in(sb_3__3__grid_top_l_in),
        .grid_right_t_in(sb_3__3__grid_right_t_in),
        .grid_right_b_in(sb_3__3__grid_right_b_in),
        .grid_bottom_r_in(sb_3__2__grid_top_r_in),
        .grid_bottom_l_in(sb_3__2__grid_top_l_in),
        .grid_left_t_in(sb_2__3__grid_right_t_in),
        .grid_left_b_in(sb_2__3__grid_right_b_in),
        .bl({bl[14204], bl[14205], bl[14206], bl[14207], bl[14208], bl[14209], bl[14210], bl[14211], bl[14212], bl[14213], bl[14214], bl[14215], bl[14216], bl[14217], bl[14218], bl[14219], bl[14220], bl[14221], bl[14222], bl[14223], bl[14224], bl[14225], bl[14226], bl[14227], bl[14228], bl[14229], bl[14230], bl[14231], bl[14232], bl[14233], bl[14234], bl[14235], bl[14236], bl[14237], bl[14238], bl[14239], bl[14240], bl[14241], bl[14242], bl[14243], bl[14244], bl[14245], bl[14246], bl[14247], bl[14248], bl[14249], bl[14250], bl[14251], bl[14252], bl[14253], bl[14254], bl[14255], bl[14256], bl[14257], bl[14258], bl[14259], bl[14260], bl[14261], bl[14262], bl[14263], bl[14264], bl[14265], bl[14266], bl[14267], bl[14268], bl[14269], bl[14270], bl[14271], bl[14272], bl[14273], bl[14274], bl[14275], bl[14276], bl[14277], bl[14278], bl[14279], bl[14280], bl[14281], bl[14282], bl[14283], bl[14284], bl[14285], bl[14286], bl[14287], bl[14288], bl[14289], bl[14290], bl[14291], bl[14292], bl[14293], bl[14294], bl[14295], bl[14296], bl[14297], bl[14298], bl[14299], bl[14300], bl[14301], bl[14302], bl[14303], bl[14304], bl[14305], bl[14306], bl[14307], bl[14308], bl[14309], bl[14310], bl[14311], bl[14312], bl[14313], bl[14314], bl[14315], bl[14316], bl[14317], bl[14318], bl[14319], bl[14320], bl[14321], bl[14322], bl[14323], bl[14324], bl[14325], bl[14326], bl[14327], bl[14328], bl[14329], bl[14330], bl[14331], bl[14332], bl[14333], bl[14334], bl[14335], bl[14336], bl[14337], bl[14338], bl[14339], bl[14340], bl[14341], bl[14342], bl[14343], bl[14344], bl[14345], bl[14346], bl[14347], bl[14348], bl[14349], bl[14350], bl[14351], bl[14352], bl[14353], bl[14354], bl[14355], bl[14356], bl[14357], bl[14358], bl[14359], bl[14360], bl[14361], bl[14362], bl[14363], bl[14364], bl[14365], bl[14366], bl[14367], bl[14368], bl[14369], bl[14370], bl[14371], bl[14372], bl[14373], bl[14374], bl[14375], bl[14376], bl[14377], bl[14378], bl[14379], bl[14380], bl[14381], bl[14382], bl[14383], bl[14384], bl[14385], bl[14386], bl[14387], bl[14388], bl[14389], bl[14390], bl[14391], bl[14392], bl[14393], bl[14394], bl[14395], bl[14396], bl[14397], bl[14398], bl[14399], bl[14400], bl[14401], bl[14402], bl[14403], bl[14404], bl[14405], bl[14406], bl[14407], bl[14408], bl[14409], bl[14410], bl[14411], bl[14412], bl[14413], bl[14414], bl[14415], bl[14416], bl[14417], bl[14418], bl[14419], bl[14420], bl[14421], bl[14422], bl[14423], bl[14424], bl[14425], bl[14426], bl[14427], bl[14428], bl[14429], bl[14430], bl[14431], bl[14432], bl[14433], bl[14434], bl[14435], bl[14436], bl[14437], bl[14438], bl[14439], bl[14440], bl[14441], bl[14442], bl[14443], bl[14444], bl[14445], bl[14446], bl[14447], bl[14448], bl[14449], bl[14450], bl[14451], bl[14452], bl[14453], bl[14454], bl[14455], bl[14456], bl[14457], bl[14458], bl[14459], bl[14460], bl[14461], bl[14462], bl[14463], bl[14464], bl[14465], bl[14466], bl[14467], bl[14468], bl[14469], bl[14470], bl[14471], bl[14472], bl[14473], bl[14474], bl[14475], bl[14476], bl[14477], bl[14478], bl[14479], bl[14480], bl[14481], bl[14482], bl[14483], bl[14484], bl[14485], bl[14486], bl[14487], bl[14488], bl[14489], bl[14490], bl[14491], bl[14492], bl[14493], bl[14494], bl[14495], bl[14496], bl[14497], bl[14498], bl[14499], bl[14500], bl[14501], bl[14502], bl[14503], bl[14504], bl[14505], bl[14506], bl[14507], bl[14508], bl[14509], bl[14510], bl[14511], bl[14512], bl[14513], bl[14514], bl[14515], bl[14516], bl[14517], bl[14518], bl[14519], bl[14520], bl[14521], bl[14522], bl[14523], bl[14524], bl[14525], bl[14526], bl[14527], bl[14528], bl[14529], bl[14530], bl[14531], bl[14532], bl[14533], bl[14534], bl[14535], bl[14536], bl[14537], bl[14538], bl[14539], bl[14540], bl[14541], bl[14542], bl[14543], bl[14544], bl[14545], bl[14546], bl[14547], bl[14548], bl[14549], bl[14550], bl[14551], bl[14552], bl[14553], bl[14554], bl[14555], bl[14556], bl[14557], bl[14558], bl[14559], bl[14560], bl[14561], bl[14562], bl[14563], bl[14564], bl[14565], bl[14566], bl[14567], bl[14568], bl[14569], bl[14570], bl[14571], bl[14572], bl[14573], bl[14574], bl[14575], bl[14576], bl[14577], bl[14578], bl[14579], bl[14580], bl[14581], bl[14582], bl[14583], bl[14584], bl[14585], bl[14586], bl[14587], bl[14588], bl[14589], bl[14590], bl[14591], bl[14592], bl[14593], bl[14594], bl[14595], bl[14596], bl[14597], bl[14598], bl[14599], bl[14600], bl[14601], bl[14602], bl[14603], bl[14604], bl[14605], bl[14606], bl[14607], bl[14608], bl[14609], bl[14610], bl[14611], bl[14612], bl[14613], bl[14614], bl[14615], bl[14616], bl[14617], bl[14618], bl[14619], bl[14620], bl[14621], bl[14622], bl[14623], bl[14624], bl[14625], bl[14626], bl[14627], bl[14628], bl[14629], bl[14630], bl[14631], bl[14632], bl[14633], bl[14634], bl[14635], bl[14636], bl[14637], bl[14638], bl[14639], bl[14640], bl[14641], bl[14642], bl[14643], bl[14644], bl[14645], bl[14646], bl[14647], bl[14648], bl[14649], bl[14650], bl[14651], bl[14652], bl[14653], bl[14654], bl[14655], bl[14656], bl[14657], bl[14658], bl[14659], bl[14660], bl[14661], bl[14662], bl[14663], bl[14664], bl[14665], bl[14666], bl[14667], bl[14668], bl[14669], bl[14670], bl[14671], bl[14672], bl[14673], bl[14674], bl[14675], bl[14676], bl[14677], bl[14678], bl[14679], bl[14680], bl[14681], bl[14682], bl[14683], bl[14684], bl[14685], bl[14686], bl[14687], bl[14688], bl[14689], bl[14690], bl[14691], bl[14692], bl[14693], bl[14694], bl[14695], bl[14696], bl[14697], bl[14698], bl[14699], bl[14700], bl[14701], bl[14702], bl[14703], bl[14704], bl[14705], bl[14706], bl[14707], bl[14708], bl[14709], bl[14710], bl[14711], bl[14712], bl[14713], bl[14714], bl[14715], bl[14716], bl[14717], bl[14718], bl[14719], bl[14720], bl[14721], bl[14722], bl[14723], bl[14724], bl[14725], bl[14726], bl[14727], bl[14728], bl[14729], bl[14730], bl[14731], bl[14732], bl[14733], bl[14734], bl[14735], bl[14736], bl[14737], bl[14738], bl[14739], bl[14740], bl[14741], bl[14742], bl[14743], bl[14744], bl[14745], bl[14746], bl[14747], bl[14748], bl[14749], bl[14750], bl[14751], bl[14752], bl[14753], bl[14754], bl[14755], bl[14756], bl[14757], bl[14758], bl[14759], bl[14760], bl[14761], bl[14762], bl[14763], bl[14764], bl[14765], bl[14766], bl[14767], bl[14768], bl[14769], bl[14770], bl[14771], bl[14772], bl[14773], bl[14774], bl[14775], bl[14776], bl[14777], bl[14778], bl[14779], bl[14780], bl[14781], bl[14782], bl[14783], bl[14784], bl[14785], bl[14786], bl[14787], bl[14788], bl[14789], bl[14790], bl[14791], bl[14792], bl[14793], bl[14794], bl[14795], bl[14796], bl[14797], bl[14798], bl[14799], bl[14800], bl[14801], bl[14802], bl[14803], bl[14804], bl[14805], bl[14806], bl[14807], bl[14808], bl[14809], bl[14810], bl[14811], bl[14812], bl[14813], bl[14814], bl[14815], bl[14816], bl[14817], bl[14818], bl[14819], bl[14820], bl[14821], bl[14822], bl[14823], bl[14824], bl[14825], bl[14826], bl[14827], bl[14828], bl[14829], bl[14830], bl[14831], bl[14832], bl[14833], bl[14834], bl[14835], bl[14836], bl[14837], bl[14838], bl[14839], bl[14840], bl[14841], bl[14842], bl[14843], bl[14844], bl[14845], bl[14846], bl[14847], bl[14848], bl[14849], bl[14850], bl[14851], bl[14852], bl[14853], bl[14854], bl[14855], bl[14856], bl[14857], bl[14858], bl[14859], bl[14860], bl[14861], bl[14862], bl[14863], bl[14864], bl[14865], bl[14866], bl[14867], bl[14868], bl[14869], bl[14870], bl[14871], bl[14872], bl[14873], bl[14874], bl[14875], bl[14876], bl[14877], bl[14878], bl[14879], bl[14880], bl[14881], bl[14882], bl[14883], bl[14884], bl[14885], bl[14886], bl[14887], bl[14888], bl[14889], bl[14890], bl[14891], bl[14892], bl[14893], bl[14894], bl[14895], bl[14896], bl[14897], bl[14898], bl[14899], bl[14900], bl[14901], bl[14902], bl[14903], bl[14904], bl[14905], bl[14906], bl[14907], bl[14908], bl[14909], bl[14910], bl[14911], bl[14912], bl[14913], bl[14914], bl[14915], bl[14916], bl[14917], bl[14918], bl[14919], bl[14920], bl[14921], bl[14922], bl[14923], bl[14924], bl[14925], bl[14926], bl[14927], bl[14928], bl[14929], bl[14930], bl[14931], bl[14932], bl[14933], bl[14934], bl[14935], bl[14936], bl[14937], bl[14938], bl[14939], bl[14940], bl[14941], bl[14942], bl[14943], bl[14944], bl[14945], bl[14946], bl[14947], bl[14948], bl[14949], bl[14950], bl[14951], bl[14952], bl[14953], bl[14954], bl[14955], bl[14956], bl[14957], bl[14958], bl[14959], bl[14960], bl[14961], bl[14962], bl[14963], bl[14964], bl[14965], bl[14966], bl[14967], bl[14968], bl[14969], bl[14970], bl[14971], bl[14972], bl[14973], bl[14974], bl[14975], bl[14976], bl[14977], bl[14978], bl[14979], bl[14980], bl[14981], bl[14982], bl[14983], bl[14984], bl[14985], bl[14986], bl[14987], bl[14988], bl[14989], bl[14990], bl[14991], bl[14992], bl[14993], bl[14994], bl[14995], bl[14996], bl[14997], bl[14998], bl[14999], bl[15000], bl[15001], bl[15002], bl[15003], bl[15004], bl[15005], bl[15006], bl[15007], bl[15008], bl[15009], bl[15010], bl[15011], bl[15012], bl[15013], bl[15014], bl[15015], bl[15016], bl[15017], bl[15018], bl[15019], bl[15020], bl[15021], bl[15022], bl[15023], bl[15024], bl[15025], bl[15026], bl[15027], bl[15028], bl[15029], bl[15030], bl[15031], bl[15032], bl[15033], bl[15034], bl[15035], bl[15036], bl[15037], bl[15038], bl[15039], bl[15040], bl[15041], bl[15042], bl[15043], bl[15044], bl[15045], bl[15046], bl[15047], bl[15048], bl[15049], bl[15050], bl[15051], bl[15052], bl[15053], bl[15054], bl[15055], bl[15056], bl[15057], bl[15058], bl[15059], bl[15060], bl[15061], bl[15062], bl[15063], bl[15064], bl[15065], bl[15066], bl[15067], bl[15068], bl[15069], bl[15070], bl[15071], bl[15072], bl[15073], bl[15074], bl[15075], bl[15076], bl[15077], bl[15078], bl[15079], bl[15080], bl[15081], bl[15082], bl[15083], bl[15084], bl[15085], bl[15086], bl[15087], bl[15088], bl[15089], bl[15090], bl[15091], bl[15092], bl[15093], bl[15094], bl[15095], bl[15096], bl[15097], bl[15098], bl[15099], bl[15100], bl[15101], bl[15102], bl[15103], bl[15104], bl[15105], bl[15106], bl[15107], bl[15108], bl[15109], bl[15110], bl[15111], bl[15112], bl[15113], bl[15114], bl[15115], bl[15116], bl[15117], bl[15118], bl[15119], bl[15120], bl[15121], bl[15122], bl[15123], bl[15124], bl[15125], bl[15126], bl[15127], bl[15128], bl[15129], bl[15130], bl[15131], bl[15132], bl[15133], bl[15134], bl[15135], bl[15136], bl[15137], bl[15138], bl[15139], bl[15140], bl[15141], bl[15142], bl[15143], bl[15144], bl[15145], bl[15146], bl[15147], bl[15148], bl[15149], bl[15150], bl[15151], bl[15152], bl[15153], bl[15154], bl[15155], bl[15156], bl[15157], bl[15158], bl[15159], bl[15160], bl[15161], bl[15162], bl[15163], bl[15164], bl[15165], bl[15166], bl[15167], bl[15168], bl[15169], bl[15170], bl[15171], bl[15172], bl[15173], bl[15174], bl[15175], bl[15176], bl[15177], bl[15178], bl[15179], bl[15180], bl[15181], bl[15182], bl[15183], bl[15184], bl[15185], bl[15186], bl[15187], bl[15188], bl[15189], bl[15190], bl[15191], bl[15192], bl[15193], bl[15194], bl[15195], bl[15196], bl[15197], bl[15198], bl[15199], bl[15200], bl[15201], bl[15202], bl[15203], bl[15204], bl[15205], bl[15206], bl[15207], bl[15208], bl[15209], bl[15210], bl[15211], bl[15212], bl[15213], bl[15214], bl[15215], bl[15216], bl[15217], bl[15218], bl[15219], bl[15220], bl[15221], bl[15222], bl[15223], bl[17808], bl[17809], bl[17810], bl[17811], bl[17812], bl[17813], bl[17814], bl[17815], bl[17816], bl[17817], bl[17818], bl[17819], bl[17820], bl[17821], bl[17822], bl[17823], bl[17824], bl[17825], bl[17826], bl[17827], bl[17828], bl[17829], bl[17830], bl[17831], bl[17832], bl[17833], bl[17834], bl[17835], bl[17836], bl[17837], bl[17838], bl[17839], bl[17840], bl[17841], bl[17842], bl[17843], bl[17844], bl[17845], bl[17846], bl[17847], bl[17848], bl[17849], bl[17850], bl[17851], bl[17852], bl[17853], bl[17854], bl[17855], bl[17856], bl[17857], bl[17858], bl[17859], bl[17860], bl[17861], bl[17862], bl[17863], bl[17864], bl[17865], bl[17866], bl[17867], bl[17868], bl[17869], bl[17870], bl[17871], bl[17872], bl[17873], bl[17874], bl[17875], bl[17876], bl[17877], bl[17878], bl[17879], bl[17880], bl[17881], bl[17882], bl[17883], bl[17884], bl[17885], bl[17886], bl[17887], bl[14124], bl[14125], bl[14126], bl[14127], bl[14128], bl[14129], bl[14130], bl[14131], bl[14132], bl[14133], bl[14134], bl[14135], bl[14136], bl[14137], bl[14138], bl[14139], bl[14140], bl[14141], bl[14142], bl[14143], bl[14144], bl[14145], bl[14146], bl[14147], bl[14148], bl[14149], bl[14150], bl[14151], bl[14152], bl[14153], bl[14154], bl[14155], bl[14156], bl[14157], bl[14158], bl[14159], bl[14160], bl[14161], bl[14162], bl[14163], bl[14164], bl[14165], bl[14166], bl[14167], bl[14168], bl[14169], bl[14170], bl[14171], bl[14172], bl[14173], bl[14174], bl[14175], bl[14176], bl[14177], bl[14178], bl[14179], bl[14180], bl[14181], bl[14182], bl[14183], bl[14184], bl[14185], bl[14186], bl[14187], bl[14188], bl[14189], bl[14190], bl[14191], bl[14192], bl[14193], bl[14194], bl[14195], bl[14196], bl[14197], bl[14198], bl[14199], bl[14200], bl[14201], bl[14202], bl[14203], bl[17728], bl[17729], bl[17730], bl[17731], bl[17732], bl[17733], bl[17734], bl[17735], bl[17736], bl[17737], bl[17738], bl[17739], bl[17740], bl[17741], bl[17742], bl[17743], bl[17744], bl[17745], bl[17746], bl[17747], bl[17748], bl[17749], bl[17750], bl[17751], bl[17752], bl[17753], bl[17754], bl[17755], bl[17756], bl[17757], bl[17758], bl[17759], bl[17760], bl[17761], bl[17762], bl[17763], bl[17764], bl[17765], bl[17766], bl[17767], bl[17768], bl[17769], bl[17770], bl[17771], bl[17772], bl[17773], bl[17774], bl[17775], bl[17776], bl[17777], bl[17778], bl[17779], bl[17780], bl[17781], bl[17782], bl[17783], bl[17784], bl[17785], bl[17786], bl[17787], bl[17788], bl[17789], bl[17790], bl[17791], bl[17792], bl[17793], bl[17794], bl[17795], bl[17796], bl[17797], bl[17798], bl[17799], bl[17800], bl[17801], bl[17802], bl[17803], bl[17804], bl[17805], bl[17806], bl[17807]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    right_tile tile_5__2_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_3__1__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_3__1__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_3__1__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_4__0__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_4__0__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_4__0__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_3__0__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_3__0__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_3__0__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_3__0__grid_top_r_in[1]),
        .grid_left_in(grid_clb_4__1__grid_left_in),
        .grid_bottom_in(grid_clb_4__1__grid_bottom_in),
        .chanx_left_in(sb_1__1__6_chanx_right_out),
        .chanx_left_out(cbx_1__1__9_chanx_left_out),
        .grid_top_out(grid_clb_4__2__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[56:63]),
        .io_left_in(grid_io_right_5__1__io_left_in),
        .chany_bottom_in(sb_4__0__0_chany_top_out),
        .chany_bottom_out(cby_4__1__0_chany_bottom_out),
        .chany_top_in_0(cby_4__1__1_chany_bottom_out),
        .chany_top_out_0(sb_4__1__0_chany_top_out),
        .grid_top_r_inpad(grid_io_right_5__2__io_left_in),
        .grid_top_l_in(sb_4__1__grid_top_l_in),
        .grid_bottom_l_in(sb_4__0__grid_top_l_in),
        .grid_left_t_in(sb_3__1__grid_right_t_in),
        .grid_left_b_in(sb_3__1__grid_right_b_in),
        .bl({bl[5392], bl[5393], bl[5394], bl[5395], bl[5396], bl[5397], bl[5398], bl[5399], bl[5400], bl[5401], bl[5402], bl[5403], bl[5404], bl[5405], bl[5406], bl[5407], bl[5408], bl[5409], bl[5410], bl[5411], bl[5412], bl[5413], bl[5414], bl[5415], bl[5416], bl[5417], bl[5418], bl[5419], bl[5420], bl[5421], bl[5422], bl[5423], bl[5424], bl[5425], bl[5426], bl[5427], bl[5428], bl[5429], bl[5430], bl[5431], bl[5432], bl[5433], bl[5434], bl[5435], bl[5436], bl[5437], bl[5438], bl[5439], bl[5440], bl[5441], bl[5442], bl[5443], bl[5444], bl[5445], bl[5446], bl[5447], bl[5448], bl[5449], bl[5450], bl[5451], bl[5452], bl[5453], bl[5454], bl[5455], bl[5456], bl[5457], bl[5458], bl[5459], bl[5460], bl[5461], bl[5462], bl[5463], bl[5464], bl[5465], bl[5466], bl[5467], bl[5468], bl[5469], bl[5470], bl[5471], bl[5472], bl[5473], bl[5474], bl[5475], bl[5476], bl[5477], bl[5478], bl[5479], bl[5480], bl[5481], bl[5482], bl[5483], bl[5484], bl[5485], bl[5486], bl[5487], bl[5488], bl[5489], bl[5490], bl[5491], bl[5492], bl[5493], bl[5494], bl[5495], bl[5496], bl[5497], bl[5498], bl[5499], bl[5500], bl[5501], bl[5502], bl[5503], bl[5504], bl[5505], bl[5506], bl[5507], bl[5508], bl[5509], bl[5510], bl[5511], bl[5512], bl[5513], bl[5514], bl[5515], bl[5516], bl[5517], bl[5518], bl[5519], bl[5520], bl[5521], bl[5522], bl[5523], bl[5524], bl[5525], bl[5526], bl[5527], bl[5528], bl[5529], bl[5530], bl[5531], bl[5532], bl[5533], bl[5534], bl[5535], bl[5536], bl[5537], bl[5538], bl[5539], bl[5540], bl[5541], bl[5542], bl[5543], bl[5544], bl[5545], bl[5546], bl[5547], bl[5548], bl[5549], bl[5550], bl[5551], bl[5552], bl[5553], bl[5554], bl[5555], bl[5556], bl[5557], bl[5558], bl[5559], bl[5560], bl[5561], bl[5562], bl[5563], bl[5564], bl[5565], bl[5566], bl[5567], bl[5568], bl[5569], bl[5570], bl[5571], bl[5572], bl[5573], bl[5574], bl[5575], bl[5576], bl[5577], bl[5578], bl[5579], bl[5580], bl[5581], bl[5582], bl[5583], bl[5584], bl[5585], bl[5586], bl[5587], bl[5588], bl[5589], bl[5590], bl[5591], bl[5592], bl[5593], bl[5594], bl[5595], bl[5596], bl[5597], bl[5598], bl[5599], bl[5600], bl[5601], bl[5602], bl[5603], bl[5604], bl[5605], bl[5606], bl[5607], bl[5608], bl[5609], bl[5610], bl[5611], bl[5612], bl[5613], bl[5614], bl[5615], bl[5616], bl[5617], bl[5618], bl[5619], bl[5620], bl[5621], bl[5622], bl[5623], bl[5624], bl[5625], bl[5626], bl[5627], bl[5628], bl[5629], bl[5630], bl[5631], bl[5632], bl[5633], bl[5634], bl[5635], bl[5636], bl[5637], bl[5638], bl[5639], bl[5640], bl[5641], bl[5642], bl[5643], bl[5644], bl[5645], bl[5646], bl[5647], bl[5648], bl[5649], bl[5650], bl[5651], bl[5652], bl[5653], bl[5654], bl[5655], bl[5656], bl[5657], bl[5658], bl[5659], bl[5660], bl[5661], bl[5662], bl[5663], bl[5664], bl[5665], bl[5666], bl[5667], bl[5668], bl[5669], bl[5670], bl[5671], bl[5672], bl[5673], bl[5674], bl[5675], bl[5676], bl[5677], bl[5678], bl[5679], bl[5680], bl[5681], bl[5682], bl[5683], bl[5684], bl[5685], bl[5686], bl[5687], bl[5688], bl[5689], bl[5690], bl[5691], bl[5692], bl[5693], bl[5694], bl[5695], bl[5696], bl[5697], bl[5698], bl[5699], bl[5700], bl[5701], bl[5702], bl[5703], bl[5704], bl[5705], bl[5706], bl[5707], bl[5708], bl[5709], bl[5710], bl[5711], bl[5712], bl[5713], bl[5714], bl[5715], bl[5716], bl[5717], bl[5718], bl[5719], bl[5720], bl[5721], bl[5722], bl[5723], bl[5724], bl[5725], bl[5726], bl[5727], bl[5728], bl[5729], bl[5730], bl[5731], bl[5732], bl[5733], bl[5734], bl[5735], bl[5736], bl[5737], bl[5738], bl[5739], bl[5740], bl[5741], bl[5742], bl[5743], bl[5744], bl[5745], bl[5746], bl[5747], bl[5748], bl[5749], bl[5750], bl[5751], bl[5752], bl[5753], bl[5754], bl[5755], bl[5756], bl[5757], bl[5758], bl[5759], bl[5760], bl[5761], bl[5762], bl[5763], bl[5764], bl[5765], bl[5766], bl[5767], bl[5768], bl[5769], bl[5770], bl[5771], bl[5772], bl[5773], bl[5774], bl[5775], bl[5776], bl[5777], bl[5778], bl[5779], bl[5780], bl[5781], bl[5782], bl[5783], bl[5784], bl[5785], bl[5786], bl[5787], bl[5788], bl[5789], bl[5790], bl[5791], bl[5792], bl[5793], bl[5794], bl[5795], bl[5796], bl[5797], bl[5798], bl[5799], bl[5800], bl[5801], bl[5802], bl[5803], bl[5804], bl[5805], bl[5806], bl[5807], bl[5808], bl[5809], bl[5810], bl[5811], bl[5812], bl[5813], bl[5814], bl[5815], bl[5816], bl[5817], bl[5818], bl[5819], bl[5820], bl[5821], bl[5822], bl[5823], bl[5824], bl[5825], bl[5826], bl[5827], bl[5828], bl[5829], bl[5830], bl[5831], bl[5832], bl[5833], bl[5834], bl[5835], bl[5836], bl[5837], bl[5838], bl[5839], bl[5840], bl[5841], bl[5842], bl[5843], bl[5844], bl[5845], bl[5846], bl[5847], bl[5848], bl[5849], bl[5850], bl[5851], bl[5852], bl[5853], bl[5854], bl[5855], bl[5856], bl[5857], bl[5858], bl[5859], bl[5860], bl[5861], bl[5862], bl[5863], bl[5864], bl[5865], bl[5866], bl[5867], bl[5868], bl[5869], bl[5870], bl[5871], bl[5872], bl[5873], bl[5874], bl[5875], bl[5876], bl[5877], bl[5878], bl[5879], bl[5880], bl[5881], bl[5882], bl[5883], bl[5884], bl[5885], bl[5886], bl[5887], bl[5888], bl[5889], bl[5890], bl[5891], bl[5892], bl[5893], bl[5894], bl[5895], bl[5896], bl[5897], bl[5898], bl[5899], bl[5900], bl[5901], bl[5902], bl[5903], bl[5904], bl[5905], bl[5906], bl[5907], bl[5908], bl[5909], bl[5910], bl[5911], bl[5912], bl[5913], bl[5914], bl[5915], bl[5916], bl[5917], bl[5918], bl[5919], bl[5920], bl[5921], bl[5922], bl[5923], bl[5924], bl[5925], bl[5926], bl[5927], bl[5928], bl[5929], bl[5930], bl[5931], bl[5932], bl[5933], bl[5934], bl[5935], bl[5936], bl[5937], bl[5938], bl[5939], bl[5940], bl[5941], bl[5942], bl[5943], bl[5944], bl[5945], bl[5946], bl[5947], bl[5948], bl[5949], bl[5950], bl[5951], bl[5952], bl[5953], bl[5954], bl[5955], bl[5956], bl[5957], bl[5958], bl[5959], bl[5960], bl[5961], bl[5962], bl[5963], bl[5964], bl[5965], bl[5966], bl[5967], bl[5968], bl[5969], bl[5970], bl[5971], bl[5972], bl[5973], bl[5974], bl[5975], bl[5976], bl[5977], bl[5978], bl[5979], bl[5980], bl[5981], bl[5982], bl[5983], bl[5984], bl[5985], bl[5986], bl[5987], bl[5988], bl[5989], bl[5990], bl[5991], bl[5992], bl[5993], bl[5994], bl[5995], bl[5996], bl[5997], bl[5998], bl[5999], bl[6000], bl[6001], bl[6002], bl[6003], bl[6004], bl[6005], bl[6006], bl[6007], bl[6008], bl[6009], bl[6010], bl[6011], bl[6012], bl[6013], bl[6014], bl[6015], bl[6016], bl[6017], bl[6018], bl[6019], bl[6020], bl[6021], bl[6022], bl[6023], bl[6024], bl[6025], bl[6026], bl[6027], bl[6028], bl[6029], bl[6030], bl[6031], bl[6032], bl[6033], bl[6034], bl[6035], bl[6036], bl[6037], bl[6038], bl[6039], bl[6040], bl[6041], bl[6042], bl[6043], bl[6044], bl[6045], bl[6046], bl[6047], bl[6048], bl[6049], bl[6050], bl[6051], bl[6052], bl[6053], bl[6054], bl[6055], bl[6056], bl[6057], bl[6058], bl[6059], bl[6060], bl[6061], bl[6062], bl[6063], bl[6064], bl[6065], bl[6066], bl[6067], bl[6068], bl[6069], bl[6070], bl[6071], bl[6072], bl[6073], bl[6074], bl[6075], bl[6076], bl[6077], bl[6078], bl[6079], bl[6080], bl[6081], bl[6082], bl[6083], bl[6084], bl[6085], bl[6086], bl[6087], bl[6088], bl[6089], bl[6090], bl[6091], bl[6092], bl[6093], bl[6094], bl[6095], bl[6096], bl[6097], bl[6098], bl[6099], bl[6100], bl[6101], bl[6102], bl[6103], bl[6104], bl[6105], bl[6106], bl[6107], bl[6108], bl[6109], bl[6110], bl[6111], bl[6112], bl[6113], bl[6114], bl[6115], bl[6116], bl[6117], bl[6118], bl[6119], bl[6120], bl[6121], bl[6122], bl[6123], bl[6124], bl[6125], bl[6126], bl[6127], bl[6128], bl[6129], bl[6130], bl[6131], bl[6132], bl[6133], bl[6134], bl[6135], bl[6136], bl[6137], bl[6138], bl[6139], bl[6140], bl[6141], bl[6142], bl[6143], bl[6144], bl[6145], bl[6146], bl[6147], bl[6148], bl[6149], bl[6150], bl[6151], bl[6152], bl[6153], bl[6154], bl[6155], bl[6156], bl[6157], bl[6158], bl[6159], bl[6160], bl[6161], bl[6162], bl[6163], bl[6164], bl[6165], bl[6166], bl[6167], bl[6168], bl[6169], bl[6170], bl[6171], bl[6172], bl[6173], bl[6174], bl[6175], bl[6176], bl[6177], bl[6178], bl[6179], bl[6180], bl[6181], bl[6182], bl[6183], bl[6184], bl[6185], bl[6186], bl[6187], bl[6188], bl[6189], bl[6190], bl[6191], bl[6192], bl[6193], bl[6194], bl[6195], bl[6196], bl[6197], bl[6198], bl[6199], bl[6200], bl[6201], bl[6202], bl[6203], bl[6204], bl[6205], bl[6206], bl[6207], bl[6208], bl[6209], bl[6210], bl[6211], bl[6212], bl[6213], bl[6214], bl[6215], bl[6216], bl[6217], bl[6218], bl[6219], bl[6220], bl[6221], bl[6222], bl[6223], bl[6224], bl[6225], bl[6226], bl[6227], bl[6228], bl[6229], bl[6230], bl[6231], bl[6232], bl[6233], bl[6234], bl[6235], bl[6236], bl[6237], bl[6238], bl[6239], bl[6240], bl[6241], bl[6242], bl[6243], bl[6244], bl[6245], bl[6246], bl[6247], bl[6248], bl[6249], bl[6250], bl[6251], bl[6252], bl[6253], bl[6254], bl[6255], bl[6256], bl[6257], bl[6258], bl[6259], bl[6260], bl[6261], bl[6262], bl[6263], bl[6264], bl[6265], bl[6266], bl[6267], bl[6268], bl[6269], bl[6270], bl[6271], bl[6272], bl[6273], bl[6274], bl[6275], bl[6276], bl[6277], bl[6278], bl[6279], bl[6280], bl[6281], bl[6282], bl[6283], bl[6284], bl[6285], bl[6286], bl[6287], bl[6288], bl[6289], bl[6290], bl[6291], bl[6292], bl[6293], bl[6294], bl[6295], bl[6296], bl[6297], bl[6298], bl[6299], bl[6300], bl[6301], bl[6302], bl[6303], bl[6304], bl[6305], bl[6306], bl[6307], bl[6308], bl[6309], bl[6310], bl[6311], bl[6312], bl[6313], bl[6314], bl[6315], bl[6316], bl[6317], bl[6318], bl[6319], bl[6320], bl[6321], bl[6322], bl[6323], bl[6324], bl[6325], bl[6326], bl[6327], bl[6328], bl[6329], bl[6330], bl[6331], bl[6332], bl[6333], bl[6334], bl[6335], bl[6336], bl[6337], bl[6338], bl[6339], bl[6340], bl[6341], bl[6342], bl[6343], bl[6344], bl[6345], bl[6346], bl[6347], bl[6348], bl[6349], bl[6350], bl[6351], bl[6352], bl[6353], bl[6354], bl[6355], bl[6356], bl[6357], bl[6358], bl[6359], bl[6360], bl[6361], bl[6362], bl[6363], bl[6364], bl[6365], bl[6366], bl[6367], bl[6368], bl[6369], bl[6370], bl[6371], bl[6372], bl[6373], bl[6374], bl[6375], bl[6376], bl[6377], bl[6378], bl[6379], bl[6380], bl[6381], bl[6382], bl[6383], bl[6384], bl[6385], bl[6386], bl[6387], bl[6388], bl[6389], bl[6390], bl[6391], bl[6392], bl[6393], bl[6394], bl[6395], bl[6396], bl[6397], bl[6398], bl[6399], bl[6400], bl[6401], bl[6402], bl[6403], bl[6404], bl[6405], bl[6406], bl[6407], bl[6408], bl[6409], bl[6410], bl[6411], bl[6492], bl[6493], bl[6494], bl[6495], bl[6496], bl[6497], bl[6498], bl[6499], bl[6500], bl[6501], bl[6502], bl[6503], bl[6504], bl[6505], bl[6506], bl[6507], bl[6508], bl[6509], bl[6510], bl[6511], bl[6512], bl[6513], bl[6514], bl[6515], bl[6516], bl[6517], bl[6518], bl[6519], bl[6520], bl[6521], bl[6522], bl[6523], bl[6524], bl[6525], bl[6526], bl[6527], bl[6528], bl[6529], bl[6530], bl[6531], bl[6532], bl[6533], bl[6534], bl[6535], bl[6536], bl[6537], bl[6538], bl[6539], bl[6540], bl[6541], bl[6542], bl[6543], bl[6544], bl[6545], bl[6546], bl[6547], bl[6548], bl[6549], bl[6550], bl[6551], bl[6552], bl[6553], bl[6554], bl[6555], bl[6556], bl[6557], bl[6558], bl[6559], bl[6560], bl[6561], bl[6562], bl[6563], bl[6564], bl[6565], bl[6566], bl[6567], bl[6568], bl[6569], bl[6570], bl[6571], bl[32], bl[33], bl[34], bl[35], bl[36], bl[37], bl[38], bl[39], bl[5320], bl[5321], bl[5322], bl[5323], bl[5324], bl[5325], bl[5326], bl[5327], bl[5328], bl[5329], bl[5330], bl[5331], bl[5332], bl[5333], bl[5334], bl[5335], bl[5336], bl[5337], bl[5338], bl[5339], bl[5340], bl[5341], bl[5342], bl[5343], bl[5344], bl[5345], bl[5346], bl[5347], bl[5348], bl[5349], bl[5350], bl[5351], bl[5352], bl[5353], bl[5354], bl[5355], bl[5356], bl[5357], bl[5358], bl[5359], bl[5360], bl[5361], bl[5362], bl[5363], bl[5364], bl[5365], bl[5366], bl[5367], bl[5368], bl[5369], bl[5370], bl[5371], bl[5372], bl[5373], bl[5374], bl[5375], bl[5376], bl[5377], bl[5378], bl[5379], bl[5380], bl[5381], bl[5382], bl[5383], bl[5384], bl[5385], bl[5386], bl[5387], bl[5388], bl[5389], bl[5390], bl[5391], bl[6412], bl[6413], bl[6414], bl[6415], bl[6416], bl[6417], bl[6418], bl[6419], bl[6420], bl[6421], bl[6422], bl[6423], bl[6424], bl[6425], bl[6426], bl[6427], bl[6428], bl[6429], bl[6430], bl[6431], bl[6432], bl[6433], bl[6434], bl[6435], bl[6436], bl[6437], bl[6438], bl[6439], bl[6440], bl[6441], bl[6442], bl[6443], bl[6444], bl[6445], bl[6446], bl[6447], bl[6448], bl[6449], bl[6450], bl[6451], bl[6452], bl[6453], bl[6454], bl[6455], bl[6456], bl[6457], bl[6458], bl[6459], bl[6460], bl[6461], bl[6462], bl[6463], bl[6464], bl[6465], bl[6466], bl[6467], bl[6468], bl[6469], bl[6470], bl[6471], bl[6472], bl[6473], bl[6474], bl[6475], bl[6476], bl[6477], bl[6478], bl[6479], bl[6480], bl[6481], bl[6482], bl[6483], bl[6484], bl[6485], bl[6486], bl[6487], bl[6488], bl[6489], bl[6490], bl[6491]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    right_tile tile_5__3_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_3__2__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_3__2__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_3__2__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_4__1__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_4__1__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_4__1__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_3__1__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_3__1__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_3__1__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_3__1__grid_top_r_in[1]),
        .grid_left_in(grid_clb_4__2__grid_left_in),
        .grid_bottom_in(grid_clb_4__2__grid_bottom_in),
        .chanx_left_in(sb_1__1__7_chanx_right_out),
        .chanx_left_out(cbx_1__1__10_chanx_left_out),
        .grid_top_out(grid_clb_4__3__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[48:55]),
        .io_left_in(grid_io_right_5__2__io_left_in),
        .chany_bottom_in(sb_4__1__0_chany_top_out),
        .chany_bottom_out(cby_4__1__1_chany_bottom_out),
        .chany_top_in_0(cby_4__1__2_chany_bottom_out),
        .chany_top_out_0(sb_4__1__1_chany_top_out),
        .grid_top_r_inpad(grid_io_right_5__3__io_left_in),
        .grid_top_l_in(sb_4__2__grid_top_l_in),
        .grid_bottom_l_in(sb_4__1__grid_top_l_in),
        .grid_left_t_in(sb_3__2__grid_right_t_in),
        .grid_left_b_in(sb_3__2__grid_right_b_in),
        .bl({bl[6644], bl[6645], bl[6646], bl[6647], bl[6648], bl[6649], bl[6650], bl[6651], bl[6652], bl[6653], bl[6654], bl[6655], bl[6656], bl[6657], bl[6658], bl[6659], bl[6660], bl[6661], bl[6662], bl[6663], bl[6664], bl[6665], bl[6666], bl[6667], bl[6668], bl[6669], bl[6670], bl[6671], bl[6672], bl[6673], bl[6674], bl[6675], bl[6676], bl[6677], bl[6678], bl[6679], bl[6680], bl[6681], bl[6682], bl[6683], bl[6684], bl[6685], bl[6686], bl[6687], bl[6688], bl[6689], bl[6690], bl[6691], bl[6692], bl[6693], bl[6694], bl[6695], bl[6696], bl[6697], bl[6698], bl[6699], bl[6700], bl[6701], bl[6702], bl[6703], bl[6704], bl[6705], bl[6706], bl[6707], bl[6708], bl[6709], bl[6710], bl[6711], bl[6712], bl[6713], bl[6714], bl[6715], bl[6716], bl[6717], bl[6718], bl[6719], bl[6720], bl[6721], bl[6722], bl[6723], bl[6724], bl[6725], bl[6726], bl[6727], bl[6728], bl[6729], bl[6730], bl[6731], bl[6732], bl[6733], bl[6734], bl[6735], bl[6736], bl[6737], bl[6738], bl[6739], bl[6740], bl[6741], bl[6742], bl[6743], bl[6744], bl[6745], bl[6746], bl[6747], bl[6748], bl[6749], bl[6750], bl[6751], bl[6752], bl[6753], bl[6754], bl[6755], bl[6756], bl[6757], bl[6758], bl[6759], bl[6760], bl[6761], bl[6762], bl[6763], bl[6764], bl[6765], bl[6766], bl[6767], bl[6768], bl[6769], bl[6770], bl[6771], bl[6772], bl[6773], bl[6774], bl[6775], bl[6776], bl[6777], bl[6778], bl[6779], bl[6780], bl[6781], bl[6782], bl[6783], bl[6784], bl[6785], bl[6786], bl[6787], bl[6788], bl[6789], bl[6790], bl[6791], bl[6792], bl[6793], bl[6794], bl[6795], bl[6796], bl[6797], bl[6798], bl[6799], bl[6800], bl[6801], bl[6802], bl[6803], bl[6804], bl[6805], bl[6806], bl[6807], bl[6808], bl[6809], bl[6810], bl[6811], bl[6812], bl[6813], bl[6814], bl[6815], bl[6816], bl[6817], bl[6818], bl[6819], bl[6820], bl[6821], bl[6822], bl[6823], bl[6824], bl[6825], bl[6826], bl[6827], bl[6828], bl[6829], bl[6830], bl[6831], bl[6832], bl[6833], bl[6834], bl[6835], bl[6836], bl[6837], bl[6838], bl[6839], bl[6840], bl[6841], bl[6842], bl[6843], bl[6844], bl[6845], bl[6846], bl[6847], bl[6848], bl[6849], bl[6850], bl[6851], bl[6852], bl[6853], bl[6854], bl[6855], bl[6856], bl[6857], bl[6858], bl[6859], bl[6860], bl[6861], bl[6862], bl[6863], bl[6864], bl[6865], bl[6866], bl[6867], bl[6868], bl[6869], bl[6870], bl[6871], bl[6872], bl[6873], bl[6874], bl[6875], bl[6876], bl[6877], bl[6878], bl[6879], bl[6880], bl[6881], bl[6882], bl[6883], bl[6884], bl[6885], bl[6886], bl[6887], bl[6888], bl[6889], bl[6890], bl[6891], bl[6892], bl[6893], bl[6894], bl[6895], bl[6896], bl[6897], bl[6898], bl[6899], bl[6900], bl[6901], bl[6902], bl[6903], bl[6904], bl[6905], bl[6906], bl[6907], bl[6908], bl[6909], bl[6910], bl[6911], bl[6912], bl[6913], bl[6914], bl[6915], bl[6916], bl[6917], bl[6918], bl[6919], bl[6920], bl[6921], bl[6922], bl[6923], bl[6924], bl[6925], bl[6926], bl[6927], bl[6928], bl[6929], bl[6930], bl[6931], bl[6932], bl[6933], bl[6934], bl[6935], bl[6936], bl[6937], bl[6938], bl[6939], bl[6940], bl[6941], bl[6942], bl[6943], bl[6944], bl[6945], bl[6946], bl[6947], bl[6948], bl[6949], bl[6950], bl[6951], bl[6952], bl[6953], bl[6954], bl[6955], bl[6956], bl[6957], bl[6958], bl[6959], bl[6960], bl[6961], bl[6962], bl[6963], bl[6964], bl[6965], bl[6966], bl[6967], bl[6968], bl[6969], bl[6970], bl[6971], bl[6972], bl[6973], bl[6974], bl[6975], bl[6976], bl[6977], bl[6978], bl[6979], bl[6980], bl[6981], bl[6982], bl[6983], bl[6984], bl[6985], bl[6986], bl[6987], bl[6988], bl[6989], bl[6990], bl[6991], bl[6992], bl[6993], bl[6994], bl[6995], bl[6996], bl[6997], bl[6998], bl[6999], bl[7000], bl[7001], bl[7002], bl[7003], bl[7004], bl[7005], bl[7006], bl[7007], bl[7008], bl[7009], bl[7010], bl[7011], bl[7012], bl[7013], bl[7014], bl[7015], bl[7016], bl[7017], bl[7018], bl[7019], bl[7020], bl[7021], bl[7022], bl[7023], bl[7024], bl[7025], bl[7026], bl[7027], bl[7028], bl[7029], bl[7030], bl[7031], bl[7032], bl[7033], bl[7034], bl[7035], bl[7036], bl[7037], bl[7038], bl[7039], bl[7040], bl[7041], bl[7042], bl[7043], bl[7044], bl[7045], bl[7046], bl[7047], bl[7048], bl[7049], bl[7050], bl[7051], bl[7052], bl[7053], bl[7054], bl[7055], bl[7056], bl[7057], bl[7058], bl[7059], bl[7060], bl[7061], bl[7062], bl[7063], bl[7064], bl[7065], bl[7066], bl[7067], bl[7068], bl[7069], bl[7070], bl[7071], bl[7072], bl[7073], bl[7074], bl[7075], bl[7076], bl[7077], bl[7078], bl[7079], bl[7080], bl[7081], bl[7082], bl[7083], bl[7084], bl[7085], bl[7086], bl[7087], bl[7088], bl[7089], bl[7090], bl[7091], bl[7092], bl[7093], bl[7094], bl[7095], bl[7096], bl[7097], bl[7098], bl[7099], bl[7100], bl[7101], bl[7102], bl[7103], bl[7104], bl[7105], bl[7106], bl[7107], bl[7108], bl[7109], bl[7110], bl[7111], bl[7112], bl[7113], bl[7114], bl[7115], bl[7116], bl[7117], bl[7118], bl[7119], bl[7120], bl[7121], bl[7122], bl[7123], bl[7124], bl[7125], bl[7126], bl[7127], bl[7128], bl[7129], bl[7130], bl[7131], bl[7132], bl[7133], bl[7134], bl[7135], bl[7136], bl[7137], bl[7138], bl[7139], bl[7140], bl[7141], bl[7142], bl[7143], bl[7144], bl[7145], bl[7146], bl[7147], bl[7148], bl[7149], bl[7150], bl[7151], bl[7152], bl[7153], bl[7154], bl[7155], bl[7156], bl[7157], bl[7158], bl[7159], bl[7160], bl[7161], bl[7162], bl[7163], bl[7164], bl[7165], bl[7166], bl[7167], bl[7168], bl[7169], bl[7170], bl[7171], bl[7172], bl[7173], bl[7174], bl[7175], bl[7176], bl[7177], bl[7178], bl[7179], bl[7180], bl[7181], bl[7182], bl[7183], bl[7184], bl[7185], bl[7186], bl[7187], bl[7188], bl[7189], bl[7190], bl[7191], bl[7192], bl[7193], bl[7194], bl[7195], bl[7196], bl[7197], bl[7198], bl[7199], bl[7200], bl[7201], bl[7202], bl[7203], bl[7204], bl[7205], bl[7206], bl[7207], bl[7208], bl[7209], bl[7210], bl[7211], bl[7212], bl[7213], bl[7214], bl[7215], bl[7216], bl[7217], bl[7218], bl[7219], bl[7220], bl[7221], bl[7222], bl[7223], bl[7224], bl[7225], bl[7226], bl[7227], bl[7228], bl[7229], bl[7230], bl[7231], bl[7232], bl[7233], bl[7234], bl[7235], bl[7236], bl[7237], bl[7238], bl[7239], bl[7240], bl[7241], bl[7242], bl[7243], bl[7244], bl[7245], bl[7246], bl[7247], bl[7248], bl[7249], bl[7250], bl[7251], bl[7252], bl[7253], bl[7254], bl[7255], bl[7256], bl[7257], bl[7258], bl[7259], bl[7260], bl[7261], bl[7262], bl[7263], bl[7264], bl[7265], bl[7266], bl[7267], bl[7268], bl[7269], bl[7270], bl[7271], bl[7272], bl[7273], bl[7274], bl[7275], bl[7276], bl[7277], bl[7278], bl[7279], bl[7280], bl[7281], bl[7282], bl[7283], bl[7284], bl[7285], bl[7286], bl[7287], bl[7288], bl[7289], bl[7290], bl[7291], bl[7292], bl[7293], bl[7294], bl[7295], bl[7296], bl[7297], bl[7298], bl[7299], bl[7300], bl[7301], bl[7302], bl[7303], bl[7304], bl[7305], bl[7306], bl[7307], bl[7308], bl[7309], bl[7310], bl[7311], bl[7312], bl[7313], bl[7314], bl[7315], bl[7316], bl[7317], bl[7318], bl[7319], bl[7320], bl[7321], bl[7322], bl[7323], bl[7324], bl[7325], bl[7326], bl[7327], bl[7328], bl[7329], bl[7330], bl[7331], bl[7332], bl[7333], bl[7334], bl[7335], bl[7336], bl[7337], bl[7338], bl[7339], bl[7340], bl[7341], bl[7342], bl[7343], bl[7344], bl[7345], bl[7346], bl[7347], bl[7348], bl[7349], bl[7350], bl[7351], bl[7352], bl[7353], bl[7354], bl[7355], bl[7356], bl[7357], bl[7358], bl[7359], bl[7360], bl[7361], bl[7362], bl[7363], bl[7364], bl[7365], bl[7366], bl[7367], bl[7368], bl[7369], bl[7370], bl[7371], bl[7372], bl[7373], bl[7374], bl[7375], bl[7376], bl[7377], bl[7378], bl[7379], bl[7380], bl[7381], bl[7382], bl[7383], bl[7384], bl[7385], bl[7386], bl[7387], bl[7388], bl[7389], bl[7390], bl[7391], bl[7392], bl[7393], bl[7394], bl[7395], bl[7396], bl[7397], bl[7398], bl[7399], bl[7400], bl[7401], bl[7402], bl[7403], bl[7404], bl[7405], bl[7406], bl[7407], bl[7408], bl[7409], bl[7410], bl[7411], bl[7412], bl[7413], bl[7414], bl[7415], bl[7416], bl[7417], bl[7418], bl[7419], bl[7420], bl[7421], bl[7422], bl[7423], bl[7424], bl[7425], bl[7426], bl[7427], bl[7428], bl[7429], bl[7430], bl[7431], bl[7432], bl[7433], bl[7434], bl[7435], bl[7436], bl[7437], bl[7438], bl[7439], bl[7440], bl[7441], bl[7442], bl[7443], bl[7444], bl[7445], bl[7446], bl[7447], bl[7448], bl[7449], bl[7450], bl[7451], bl[7452], bl[7453], bl[7454], bl[7455], bl[7456], bl[7457], bl[7458], bl[7459], bl[7460], bl[7461], bl[7462], bl[7463], bl[7464], bl[7465], bl[7466], bl[7467], bl[7468], bl[7469], bl[7470], bl[7471], bl[7472], bl[7473], bl[7474], bl[7475], bl[7476], bl[7477], bl[7478], bl[7479], bl[7480], bl[7481], bl[7482], bl[7483], bl[7484], bl[7485], bl[7486], bl[7487], bl[7488], bl[7489], bl[7490], bl[7491], bl[7492], bl[7493], bl[7494], bl[7495], bl[7496], bl[7497], bl[7498], bl[7499], bl[7500], bl[7501], bl[7502], bl[7503], bl[7504], bl[7505], bl[7506], bl[7507], bl[7508], bl[7509], bl[7510], bl[7511], bl[7512], bl[7513], bl[7514], bl[7515], bl[7516], bl[7517], bl[7518], bl[7519], bl[7520], bl[7521], bl[7522], bl[7523], bl[7524], bl[7525], bl[7526], bl[7527], bl[7528], bl[7529], bl[7530], bl[7531], bl[7532], bl[7533], bl[7534], bl[7535], bl[7536], bl[7537], bl[7538], bl[7539], bl[7540], bl[7541], bl[7542], bl[7543], bl[7544], bl[7545], bl[7546], bl[7547], bl[7548], bl[7549], bl[7550], bl[7551], bl[7552], bl[7553], bl[7554], bl[7555], bl[7556], bl[7557], bl[7558], bl[7559], bl[7560], bl[7561], bl[7562], bl[7563], bl[7564], bl[7565], bl[7566], bl[7567], bl[7568], bl[7569], bl[7570], bl[7571], bl[7572], bl[7573], bl[7574], bl[7575], bl[7576], bl[7577], bl[7578], bl[7579], bl[7580], bl[7581], bl[7582], bl[7583], bl[7584], bl[7585], bl[7586], bl[7587], bl[7588], bl[7589], bl[7590], bl[7591], bl[7592], bl[7593], bl[7594], bl[7595], bl[7596], bl[7597], bl[7598], bl[7599], bl[7600], bl[7601], bl[7602], bl[7603], bl[7604], bl[7605], bl[7606], bl[7607], bl[7608], bl[7609], bl[7610], bl[7611], bl[7612], bl[7613], bl[7614], bl[7615], bl[7616], bl[7617], bl[7618], bl[7619], bl[7620], bl[7621], bl[7622], bl[7623], bl[7624], bl[7625], bl[7626], bl[7627], bl[7628], bl[7629], bl[7630], bl[7631], bl[7632], bl[7633], bl[7634], bl[7635], bl[7636], bl[7637], bl[7638], bl[7639], bl[7640], bl[7641], bl[7642], bl[7643], bl[7644], bl[7645], bl[7646], bl[7647], bl[7648], bl[7649], bl[7650], bl[7651], bl[7652], bl[7653], bl[7654], bl[7655], bl[7656], bl[7657], bl[7658], bl[7659], bl[7660], bl[7661], bl[7662], bl[7663], bl[15304], bl[15305], bl[15306], bl[15307], bl[15308], bl[15309], bl[15310], bl[15311], bl[15312], bl[15313], bl[15314], bl[15315], bl[15316], bl[15317], bl[15318], bl[15319], bl[15320], bl[15321], bl[15322], bl[15323], bl[15324], bl[15325], bl[15326], bl[15327], bl[15328], bl[15329], bl[15330], bl[15331], bl[15332], bl[15333], bl[15334], bl[15335], bl[15336], bl[15337], bl[15338], bl[15339], bl[15340], bl[15341], bl[15342], bl[15343], bl[15344], bl[15345], bl[15346], bl[15347], bl[15348], bl[15349], bl[15350], bl[15351], bl[15352], bl[15353], bl[15354], bl[15355], bl[15356], bl[15357], bl[15358], bl[15359], bl[15360], bl[15361], bl[15362], bl[15363], bl[15364], bl[15365], bl[15366], bl[15367], bl[15368], bl[15369], bl[15370], bl[15371], bl[15372], bl[15373], bl[15374], bl[15375], bl[15376], bl[15377], bl[15378], bl[15379], bl[15380], bl[15381], bl[15382], bl[15383], bl[40], bl[41], bl[42], bl[43], bl[44], bl[45], bl[46], bl[47], bl[6572], bl[6573], bl[6574], bl[6575], bl[6576], bl[6577], bl[6578], bl[6579], bl[6580], bl[6581], bl[6582], bl[6583], bl[6584], bl[6585], bl[6586], bl[6587], bl[6588], bl[6589], bl[6590], bl[6591], bl[6592], bl[6593], bl[6594], bl[6595], bl[6596], bl[6597], bl[6598], bl[6599], bl[6600], bl[6601], bl[6602], bl[6603], bl[6604], bl[6605], bl[6606], bl[6607], bl[6608], bl[6609], bl[6610], bl[6611], bl[6612], bl[6613], bl[6614], bl[6615], bl[6616], bl[6617], bl[6618], bl[6619], bl[6620], bl[6621], bl[6622], bl[6623], bl[6624], bl[6625], bl[6626], bl[6627], bl[6628], bl[6629], bl[6630], bl[6631], bl[6632], bl[6633], bl[6634], bl[6635], bl[6636], bl[6637], bl[6638], bl[6639], bl[6640], bl[6641], bl[6642], bl[6643], bl[15224], bl[15225], bl[15226], bl[15227], bl[15228], bl[15229], bl[15230], bl[15231], bl[15232], bl[15233], bl[15234], bl[15235], bl[15236], bl[15237], bl[15238], bl[15239], bl[15240], bl[15241], bl[15242], bl[15243], bl[15244], bl[15245], bl[15246], bl[15247], bl[15248], bl[15249], bl[15250], bl[15251], bl[15252], bl[15253], bl[15254], bl[15255], bl[15256], bl[15257], bl[15258], bl[15259], bl[15260], bl[15261], bl[15262], bl[15263], bl[15264], bl[15265], bl[15266], bl[15267], bl[15268], bl[15269], bl[15270], bl[15271], bl[15272], bl[15273], bl[15274], bl[15275], bl[15276], bl[15277], bl[15278], bl[15279], bl[15280], bl[15281], bl[15282], bl[15283], bl[15284], bl[15285], bl[15286], bl[15287], bl[15288], bl[15289], bl[15290], bl[15291], bl[15292], bl[15293], bl[15294], bl[15295], bl[15296], bl[15297], bl[15298], bl[15299], bl[15300], bl[15301], bl[15302], bl[15303]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    right_tile tile_5__4_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_3__3__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_3__3__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_3__3__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_4__2__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_4__2__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_4__2__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_3__2__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_3__2__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_3__2__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_3__2__grid_top_r_in[1]),
        .grid_left_in(grid_clb_4__3__grid_left_in),
        .grid_bottom_in(grid_clb_4__3__grid_bottom_in),
        .chanx_left_in(sb_1__1__8_chanx_right_out),
        .chanx_left_out(cbx_1__1__11_chanx_left_out),
        .grid_top_out(grid_clb_4__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[40:47]),
        .io_left_in(grid_io_right_5__3__io_left_in),
        .chany_bottom_in(sb_4__1__1_chany_top_out),
        .chany_bottom_out(cby_4__1__2_chany_bottom_out),
        .chany_top_in_0(cby_4__1__3_chany_bottom_out),
        .chany_top_out_0(sb_4__1__2_chany_top_out),
        .grid_top_r_inpad(grid_io_right_5__4__io_left_in),
        .grid_top_l_in(sb_4__3__grid_top_l_in),
        .grid_bottom_l_in(sb_4__2__grid_top_l_in),
        .grid_left_t_in(sb_3__3__grid_right_t_in),
        .grid_left_b_in(sb_3__3__grid_right_b_in),
        .bl({bl[15456], bl[15457], bl[15458], bl[15459], bl[15460], bl[15461], bl[15462], bl[15463], bl[15464], bl[15465], bl[15466], bl[15467], bl[15468], bl[15469], bl[15470], bl[15471], bl[15472], bl[15473], bl[15474], bl[15475], bl[15476], bl[15477], bl[15478], bl[15479], bl[15480], bl[15481], bl[15482], bl[15483], bl[15484], bl[15485], bl[15486], bl[15487], bl[15488], bl[15489], bl[15490], bl[15491], bl[15492], bl[15493], bl[15494], bl[15495], bl[15496], bl[15497], bl[15498], bl[15499], bl[15500], bl[15501], bl[15502], bl[15503], bl[15504], bl[15505], bl[15506], bl[15507], bl[15508], bl[15509], bl[15510], bl[15511], bl[15512], bl[15513], bl[15514], bl[15515], bl[15516], bl[15517], bl[15518], bl[15519], bl[15520], bl[15521], bl[15522], bl[15523], bl[15524], bl[15525], bl[15526], bl[15527], bl[15528], bl[15529], bl[15530], bl[15531], bl[15532], bl[15533], bl[15534], bl[15535], bl[15536], bl[15537], bl[15538], bl[15539], bl[15540], bl[15541], bl[15542], bl[15543], bl[15544], bl[15545], bl[15546], bl[15547], bl[15548], bl[15549], bl[15550], bl[15551], bl[15552], bl[15553], bl[15554], bl[15555], bl[15556], bl[15557], bl[15558], bl[15559], bl[15560], bl[15561], bl[15562], bl[15563], bl[15564], bl[15565], bl[15566], bl[15567], bl[15568], bl[15569], bl[15570], bl[15571], bl[15572], bl[15573], bl[15574], bl[15575], bl[15576], bl[15577], bl[15578], bl[15579], bl[15580], bl[15581], bl[15582], bl[15583], bl[15584], bl[15585], bl[15586], bl[15587], bl[15588], bl[15589], bl[15590], bl[15591], bl[15592], bl[15593], bl[15594], bl[15595], bl[15596], bl[15597], bl[15598], bl[15599], bl[15600], bl[15601], bl[15602], bl[15603], bl[15604], bl[15605], bl[15606], bl[15607], bl[15608], bl[15609], bl[15610], bl[15611], bl[15612], bl[15613], bl[15614], bl[15615], bl[15616], bl[15617], bl[15618], bl[15619], bl[15620], bl[15621], bl[15622], bl[15623], bl[15624], bl[15625], bl[15626], bl[15627], bl[15628], bl[15629], bl[15630], bl[15631], bl[15632], bl[15633], bl[15634], bl[15635], bl[15636], bl[15637], bl[15638], bl[15639], bl[15640], bl[15641], bl[15642], bl[15643], bl[15644], bl[15645], bl[15646], bl[15647], bl[15648], bl[15649], bl[15650], bl[15651], bl[15652], bl[15653], bl[15654], bl[15655], bl[15656], bl[15657], bl[15658], bl[15659], bl[15660], bl[15661], bl[15662], bl[15663], bl[15664], bl[15665], bl[15666], bl[15667], bl[15668], bl[15669], bl[15670], bl[15671], bl[15672], bl[15673], bl[15674], bl[15675], bl[15676], bl[15677], bl[15678], bl[15679], bl[15680], bl[15681], bl[15682], bl[15683], bl[15684], bl[15685], bl[15686], bl[15687], bl[15688], bl[15689], bl[15690], bl[15691], bl[15692], bl[15693], bl[15694], bl[15695], bl[15696], bl[15697], bl[15698], bl[15699], bl[15700], bl[15701], bl[15702], bl[15703], bl[15704], bl[15705], bl[15706], bl[15707], bl[15708], bl[15709], bl[15710], bl[15711], bl[15712], bl[15713], bl[15714], bl[15715], bl[15716], bl[15717], bl[15718], bl[15719], bl[15720], bl[15721], bl[15722], bl[15723], bl[15724], bl[15725], bl[15726], bl[15727], bl[15728], bl[15729], bl[15730], bl[15731], bl[15732], bl[15733], bl[15734], bl[15735], bl[15736], bl[15737], bl[15738], bl[15739], bl[15740], bl[15741], bl[15742], bl[15743], bl[15744], bl[15745], bl[15746], bl[15747], bl[15748], bl[15749], bl[15750], bl[15751], bl[15752], bl[15753], bl[15754], bl[15755], bl[15756], bl[15757], bl[15758], bl[15759], bl[15760], bl[15761], bl[15762], bl[15763], bl[15764], bl[15765], bl[15766], bl[15767], bl[15768], bl[15769], bl[15770], bl[15771], bl[15772], bl[15773], bl[15774], bl[15775], bl[15776], bl[15777], bl[15778], bl[15779], bl[15780], bl[15781], bl[15782], bl[15783], bl[15784], bl[15785], bl[15786], bl[15787], bl[15788], bl[15789], bl[15790], bl[15791], bl[15792], bl[15793], bl[15794], bl[15795], bl[15796], bl[15797], bl[15798], bl[15799], bl[15800], bl[15801], bl[15802], bl[15803], bl[15804], bl[15805], bl[15806], bl[15807], bl[15808], bl[15809], bl[15810], bl[15811], bl[15812], bl[15813], bl[15814], bl[15815], bl[15816], bl[15817], bl[15818], bl[15819], bl[15820], bl[15821], bl[15822], bl[15823], bl[15824], bl[15825], bl[15826], bl[15827], bl[15828], bl[15829], bl[15830], bl[15831], bl[15832], bl[15833], bl[15834], bl[15835], bl[15836], bl[15837], bl[15838], bl[15839], bl[15840], bl[15841], bl[15842], bl[15843], bl[15844], bl[15845], bl[15846], bl[15847], bl[15848], bl[15849], bl[15850], bl[15851], bl[15852], bl[15853], bl[15854], bl[15855], bl[15856], bl[15857], bl[15858], bl[15859], bl[15860], bl[15861], bl[15862], bl[15863], bl[15864], bl[15865], bl[15866], bl[15867], bl[15868], bl[15869], bl[15870], bl[15871], bl[15872], bl[15873], bl[15874], bl[15875], bl[15876], bl[15877], bl[15878], bl[15879], bl[15880], bl[15881], bl[15882], bl[15883], bl[15884], bl[15885], bl[15886], bl[15887], bl[15888], bl[15889], bl[15890], bl[15891], bl[15892], bl[15893], bl[15894], bl[15895], bl[15896], bl[15897], bl[15898], bl[15899], bl[15900], bl[15901], bl[15902], bl[15903], bl[15904], bl[15905], bl[15906], bl[15907], bl[15908], bl[15909], bl[15910], bl[15911], bl[15912], bl[15913], bl[15914], bl[15915], bl[15916], bl[15917], bl[15918], bl[15919], bl[15920], bl[15921], bl[15922], bl[15923], bl[15924], bl[15925], bl[15926], bl[15927], bl[15928], bl[15929], bl[15930], bl[15931], bl[15932], bl[15933], bl[15934], bl[15935], bl[15936], bl[15937], bl[15938], bl[15939], bl[15940], bl[15941], bl[15942], bl[15943], bl[15944], bl[15945], bl[15946], bl[15947], bl[15948], bl[15949], bl[15950], bl[15951], bl[15952], bl[15953], bl[15954], bl[15955], bl[15956], bl[15957], bl[15958], bl[15959], bl[15960], bl[15961], bl[15962], bl[15963], bl[15964], bl[15965], bl[15966], bl[15967], bl[15968], bl[15969], bl[15970], bl[15971], bl[15972], bl[15973], bl[15974], bl[15975], bl[15976], bl[15977], bl[15978], bl[15979], bl[15980], bl[15981], bl[15982], bl[15983], bl[15984], bl[15985], bl[15986], bl[15987], bl[15988], bl[15989], bl[15990], bl[15991], bl[15992], bl[15993], bl[15994], bl[15995], bl[15996], bl[15997], bl[15998], bl[15999], bl[16000], bl[16001], bl[16002], bl[16003], bl[16004], bl[16005], bl[16006], bl[16007], bl[16008], bl[16009], bl[16010], bl[16011], bl[16012], bl[16013], bl[16014], bl[16015], bl[16016], bl[16017], bl[16018], bl[16019], bl[16020], bl[16021], bl[16022], bl[16023], bl[16024], bl[16025], bl[16026], bl[16027], bl[16028], bl[16029], bl[16030], bl[16031], bl[16032], bl[16033], bl[16034], bl[16035], bl[16036], bl[16037], bl[16038], bl[16039], bl[16040], bl[16041], bl[16042], bl[16043], bl[16044], bl[16045], bl[16046], bl[16047], bl[16048], bl[16049], bl[16050], bl[16051], bl[16052], bl[16053], bl[16054], bl[16055], bl[16056], bl[16057], bl[16058], bl[16059], bl[16060], bl[16061], bl[16062], bl[16063], bl[16064], bl[16065], bl[16066], bl[16067], bl[16068], bl[16069], bl[16070], bl[16071], bl[16072], bl[16073], bl[16074], bl[16075], bl[16076], bl[16077], bl[16078], bl[16079], bl[16080], bl[16081], bl[16082], bl[16083], bl[16084], bl[16085], bl[16086], bl[16087], bl[16088], bl[16089], bl[16090], bl[16091], bl[16092], bl[16093], bl[16094], bl[16095], bl[16096], bl[16097], bl[16098], bl[16099], bl[16100], bl[16101], bl[16102], bl[16103], bl[16104], bl[16105], bl[16106], bl[16107], bl[16108], bl[16109], bl[16110], bl[16111], bl[16112], bl[16113], bl[16114], bl[16115], bl[16116], bl[16117], bl[16118], bl[16119], bl[16120], bl[16121], bl[16122], bl[16123], bl[16124], bl[16125], bl[16126], bl[16127], bl[16128], bl[16129], bl[16130], bl[16131], bl[16132], bl[16133], bl[16134], bl[16135], bl[16136], bl[16137], bl[16138], bl[16139], bl[16140], bl[16141], bl[16142], bl[16143], bl[16144], bl[16145], bl[16146], bl[16147], bl[16148], bl[16149], bl[16150], bl[16151], bl[16152], bl[16153], bl[16154], bl[16155], bl[16156], bl[16157], bl[16158], bl[16159], bl[16160], bl[16161], bl[16162], bl[16163], bl[16164], bl[16165], bl[16166], bl[16167], bl[16168], bl[16169], bl[16170], bl[16171], bl[16172], bl[16173], bl[16174], bl[16175], bl[16176], bl[16177], bl[16178], bl[16179], bl[16180], bl[16181], bl[16182], bl[16183], bl[16184], bl[16185], bl[16186], bl[16187], bl[16188], bl[16189], bl[16190], bl[16191], bl[16192], bl[16193], bl[16194], bl[16195], bl[16196], bl[16197], bl[16198], bl[16199], bl[16200], bl[16201], bl[16202], bl[16203], bl[16204], bl[16205], bl[16206], bl[16207], bl[16208], bl[16209], bl[16210], bl[16211], bl[16212], bl[16213], bl[16214], bl[16215], bl[16216], bl[16217], bl[16218], bl[16219], bl[16220], bl[16221], bl[16222], bl[16223], bl[16224], bl[16225], bl[16226], bl[16227], bl[16228], bl[16229], bl[16230], bl[16231], bl[16232], bl[16233], bl[16234], bl[16235], bl[16236], bl[16237], bl[16238], bl[16239], bl[16240], bl[16241], bl[16242], bl[16243], bl[16244], bl[16245], bl[16246], bl[16247], bl[16248], bl[16249], bl[16250], bl[16251], bl[16252], bl[16253], bl[16254], bl[16255], bl[16256], bl[16257], bl[16258], bl[16259], bl[16260], bl[16261], bl[16262], bl[16263], bl[16264], bl[16265], bl[16266], bl[16267], bl[16268], bl[16269], bl[16270], bl[16271], bl[16272], bl[16273], bl[16274], bl[16275], bl[16276], bl[16277], bl[16278], bl[16279], bl[16280], bl[16281], bl[16282], bl[16283], bl[16284], bl[16285], bl[16286], bl[16287], bl[16288], bl[16289], bl[16290], bl[16291], bl[16292], bl[16293], bl[16294], bl[16295], bl[16296], bl[16297], bl[16298], bl[16299], bl[16300], bl[16301], bl[16302], bl[16303], bl[16304], bl[16305], bl[16306], bl[16307], bl[16308], bl[16309], bl[16310], bl[16311], bl[16312], bl[16313], bl[16314], bl[16315], bl[16316], bl[16317], bl[16318], bl[16319], bl[16320], bl[16321], bl[16322], bl[16323], bl[16324], bl[16325], bl[16326], bl[16327], bl[16328], bl[16329], bl[16330], bl[16331], bl[16332], bl[16333], bl[16334], bl[16335], bl[16336], bl[16337], bl[16338], bl[16339], bl[16340], bl[16341], bl[16342], bl[16343], bl[16344], bl[16345], bl[16346], bl[16347], bl[16348], bl[16349], bl[16350], bl[16351], bl[16352], bl[16353], bl[16354], bl[16355], bl[16356], bl[16357], bl[16358], bl[16359], bl[16360], bl[16361], bl[16362], bl[16363], bl[16364], bl[16365], bl[16366], bl[16367], bl[16368], bl[16369], bl[16370], bl[16371], bl[16372], bl[16373], bl[16374], bl[16375], bl[16376], bl[16377], bl[16378], bl[16379], bl[16380], bl[16381], bl[16382], bl[16383], bl[16384], bl[16385], bl[16386], bl[16387], bl[16388], bl[16389], bl[16390], bl[16391], bl[16392], bl[16393], bl[16394], bl[16395], bl[16396], bl[16397], bl[16398], bl[16399], bl[16400], bl[16401], bl[16402], bl[16403], bl[16404], bl[16405], bl[16406], bl[16407], bl[16408], bl[16409], bl[16410], bl[16411], bl[16412], bl[16413], bl[16414], bl[16415], bl[16416], bl[16417], bl[16418], bl[16419], bl[16420], bl[16421], bl[16422], bl[16423], bl[16424], bl[16425], bl[16426], bl[16427], bl[16428], bl[16429], bl[16430], bl[16431], bl[16432], bl[16433], bl[16434], bl[16435], bl[16436], bl[16437], bl[16438], bl[16439], bl[16440], bl[16441], bl[16442], bl[16443], bl[16444], bl[16445], bl[16446], bl[16447], bl[16448], bl[16449], bl[16450], bl[16451], bl[16452], bl[16453], bl[16454], bl[16455], bl[16456], bl[16457], bl[16458], bl[16459], bl[16460], bl[16461], bl[16462], bl[16463], bl[16464], bl[16465], bl[16466], bl[16467], bl[16468], bl[16469], bl[16470], bl[16471], bl[16472], bl[16473], bl[16474], bl[16475], bl[16556], bl[16557], bl[16558], bl[16559], bl[16560], bl[16561], bl[16562], bl[16563], bl[16564], bl[16565], bl[16566], bl[16567], bl[16568], bl[16569], bl[16570], bl[16571], bl[16572], bl[16573], bl[16574], bl[16575], bl[16576], bl[16577], bl[16578], bl[16579], bl[16580], bl[16581], bl[16582], bl[16583], bl[16584], bl[16585], bl[16586], bl[16587], bl[16588], bl[16589], bl[16590], bl[16591], bl[16592], bl[16593], bl[16594], bl[16595], bl[16596], bl[16597], bl[16598], bl[16599], bl[16600], bl[16601], bl[16602], bl[16603], bl[16604], bl[16605], bl[16606], bl[16607], bl[16608], bl[16609], bl[16610], bl[16611], bl[16612], bl[16613], bl[16614], bl[16615], bl[16616], bl[16617], bl[16618], bl[16619], bl[16620], bl[16621], bl[16622], bl[16623], bl[16624], bl[16625], bl[16626], bl[16627], bl[16628], bl[16629], bl[16630], bl[16631], bl[16632], bl[16633], bl[16634], bl[16635], bl[48], bl[49], bl[50], bl[51], bl[52], bl[53], bl[54], bl[55], bl[15384], bl[15385], bl[15386], bl[15387], bl[15388], bl[15389], bl[15390], bl[15391], bl[15392], bl[15393], bl[15394], bl[15395], bl[15396], bl[15397], bl[15398], bl[15399], bl[15400], bl[15401], bl[15402], bl[15403], bl[15404], bl[15405], bl[15406], bl[15407], bl[15408], bl[15409], bl[15410], bl[15411], bl[15412], bl[15413], bl[15414], bl[15415], bl[15416], bl[15417], bl[15418], bl[15419], bl[15420], bl[15421], bl[15422], bl[15423], bl[15424], bl[15425], bl[15426], bl[15427], bl[15428], bl[15429], bl[15430], bl[15431], bl[15432], bl[15433], bl[15434], bl[15435], bl[15436], bl[15437], bl[15438], bl[15439], bl[15440], bl[15441], bl[15442], bl[15443], bl[15444], bl[15445], bl[15446], bl[15447], bl[15448], bl[15449], bl[15450], bl[15451], bl[15452], bl[15453], bl[15454], bl[15455], bl[16476], bl[16477], bl[16478], bl[16479], bl[16480], bl[16481], bl[16482], bl[16483], bl[16484], bl[16485], bl[16486], bl[16487], bl[16488], bl[16489], bl[16490], bl[16491], bl[16492], bl[16493], bl[16494], bl[16495], bl[16496], bl[16497], bl[16498], bl[16499], bl[16500], bl[16501], bl[16502], bl[16503], bl[16504], bl[16505], bl[16506], bl[16507], bl[16508], bl[16509], bl[16510], bl[16511], bl[16512], bl[16513], bl[16514], bl[16515], bl[16516], bl[16517], bl[16518], bl[16519], bl[16520], bl[16521], bl[16522], bl[16523], bl[16524], bl[16525], bl[16526], bl[16527], bl[16528], bl[16529], bl[16530], bl[16531], bl[16532], bl[16533], bl[16534], bl[16535], bl[16536], bl[16537], bl[16538], bl[16539], bl[16540], bl[16541], bl[16542], bl[16543], bl[16544], bl[16545], bl[16546], bl[16547], bl[16548], bl[16549], bl[16550], bl[16551], bl[16552], bl[16553], bl[16554], bl[16555]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    top_tile tile_2__5_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_0__4__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_0__4__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_0__4__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_1__3__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_1__3__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_1__3__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_0__3__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_0__3__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_0__3__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_0__3__grid_top_r_in[1]),
        .grid_left_in(grid_clb_1__4__grid_left_in),
        .grid_bottom_in(grid_clb_1__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0:7]),
        .io_bottom_in(grid_io_top_1__5__io_bottom_in),
        .chanx_left_in(sb_0__4__0_chanx_right_out),
        .chanx_left_out(cbx_1__4__0_chanx_left_out),
        .chany_bottom_in(sb_1__1__2_chany_top_out),
        .chany_bottom_out(cby_1__1__3_chany_bottom_out),
        .grid_right_out(grid_clb_2__4__grid_left_in),
        .chanx_right_in_0(cbx_1__4__1_chanx_left_out),
        .chanx_right_out_0(sb_1__4__0_chanx_right_out),
        .grid_right_t_inpad(grid_io_top_2__5__io_bottom_in),
        .grid_right_b_in(sb_1__4__grid_right_b_in),
        .grid_bottom_r_in(sb_1__3__grid_top_r_in),
        .grid_bottom_l_in(sb_1__3__grid_top_l_in),
        .grid_left_b_in(sb_0__4__grid_right_b_in),
        .bl({bl[20488], bl[20489], bl[20490], bl[20491], bl[20492], bl[20493], bl[20494], bl[20495], bl[20496], bl[20497], bl[20498], bl[20499], bl[20500], bl[20501], bl[20502], bl[20503], bl[20504], bl[20505], bl[20506], bl[20507], bl[20508], bl[20509], bl[20510], bl[20511], bl[20512], bl[20513], bl[20514], bl[20515], bl[20516], bl[20517], bl[20518], bl[20519], bl[20520], bl[20521], bl[20522], bl[20523], bl[20524], bl[20525], bl[20526], bl[20527], bl[20528], bl[20529], bl[20530], bl[20531], bl[20532], bl[20533], bl[20534], bl[20535], bl[20536], bl[20537], bl[20538], bl[20539], bl[20540], bl[20541], bl[20542], bl[20543], bl[20544], bl[20545], bl[20546], bl[20547], bl[20548], bl[20549], bl[20550], bl[20551], bl[20552], bl[20553], bl[20554], bl[20555], bl[20556], bl[20557], bl[20558], bl[20559], bl[20560], bl[20561], bl[20562], bl[20563], bl[20564], bl[20565], bl[20566], bl[20567], bl[20568], bl[20569], bl[20570], bl[20571], bl[20572], bl[20573], bl[20574], bl[20575], bl[20576], bl[20577], bl[20578], bl[20579], bl[20580], bl[20581], bl[20582], bl[20583], bl[20584], bl[20585], bl[20586], bl[20587], bl[20588], bl[20589], bl[20590], bl[20591], bl[20592], bl[20593], bl[20594], bl[20595], bl[20596], bl[20597], bl[20598], bl[20599], bl[20600], bl[20601], bl[20602], bl[20603], bl[20604], bl[20605], bl[20606], bl[20607], bl[20608], bl[20609], bl[20610], bl[20611], bl[20612], bl[20613], bl[20614], bl[20615], bl[20616], bl[20617], bl[20618], bl[20619], bl[20620], bl[20621], bl[20622], bl[20623], bl[20624], bl[20625], bl[20626], bl[20627], bl[20628], bl[20629], bl[20630], bl[20631], bl[20632], bl[20633], bl[20634], bl[20635], bl[20636], bl[20637], bl[20638], bl[20639], bl[20640], bl[20641], bl[20642], bl[20643], bl[20644], bl[20645], bl[20646], bl[20647], bl[20648], bl[20649], bl[20650], bl[20651], bl[20652], bl[20653], bl[20654], bl[20655], bl[20656], bl[20657], bl[20658], bl[20659], bl[20660], bl[20661], bl[20662], bl[20663], bl[20664], bl[20665], bl[20666], bl[20667], bl[20668], bl[20669], bl[20670], bl[20671], bl[20672], bl[20673], bl[20674], bl[20675], bl[20676], bl[20677], bl[20678], bl[20679], bl[20680], bl[20681], bl[20682], bl[20683], bl[20684], bl[20685], bl[20686], bl[20687], bl[20688], bl[20689], bl[20690], bl[20691], bl[20692], bl[20693], bl[20694], bl[20695], bl[20696], bl[20697], bl[20698], bl[20699], bl[20700], bl[20701], bl[20702], bl[20703], bl[20704], bl[20705], bl[20706], bl[20707], bl[20708], bl[20709], bl[20710], bl[20711], bl[20712], bl[20713], bl[20714], bl[20715], bl[20716], bl[20717], bl[20718], bl[20719], bl[20720], bl[20721], bl[20722], bl[20723], bl[20724], bl[20725], bl[20726], bl[20727], bl[20728], bl[20729], bl[20730], bl[20731], bl[20732], bl[20733], bl[20734], bl[20735], bl[20736], bl[20737], bl[20738], bl[20739], bl[20740], bl[20741], bl[20742], bl[20743], bl[20744], bl[20745], bl[20746], bl[20747], bl[20748], bl[20749], bl[20750], bl[20751], bl[20752], bl[20753], bl[20754], bl[20755], bl[20756], bl[20757], bl[20758], bl[20759], bl[20760], bl[20761], bl[20762], bl[20763], bl[20764], bl[20765], bl[20766], bl[20767], bl[20768], bl[20769], bl[20770], bl[20771], bl[20772], bl[20773], bl[20774], bl[20775], bl[20776], bl[20777], bl[20778], bl[20779], bl[20780], bl[20781], bl[20782], bl[20783], bl[20784], bl[20785], bl[20786], bl[20787], bl[20788], bl[20789], bl[20790], bl[20791], bl[20792], bl[20793], bl[20794], bl[20795], bl[20796], bl[20797], bl[20798], bl[20799], bl[20800], bl[20801], bl[20802], bl[20803], bl[20804], bl[20805], bl[20806], bl[20807], bl[20808], bl[20809], bl[20810], bl[20811], bl[20812], bl[20813], bl[20814], bl[20815], bl[20816], bl[20817], bl[20818], bl[20819], bl[20820], bl[20821], bl[20822], bl[20823], bl[20824], bl[20825], bl[20826], bl[20827], bl[20828], bl[20829], bl[20830], bl[20831], bl[20832], bl[20833], bl[20834], bl[20835], bl[20836], bl[20837], bl[20838], bl[20839], bl[20840], bl[20841], bl[20842], bl[20843], bl[20844], bl[20845], bl[20846], bl[20847], bl[20848], bl[20849], bl[20850], bl[20851], bl[20852], bl[20853], bl[20854], bl[20855], bl[20856], bl[20857], bl[20858], bl[20859], bl[20860], bl[20861], bl[20862], bl[20863], bl[20864], bl[20865], bl[20866], bl[20867], bl[20868], bl[20869], bl[20870], bl[20871], bl[20872], bl[20873], bl[20874], bl[20875], bl[20876], bl[20877], bl[20878], bl[20879], bl[20880], bl[20881], bl[20882], bl[20883], bl[20884], bl[20885], bl[20886], bl[20887], bl[20888], bl[20889], bl[20890], bl[20891], bl[20892], bl[20893], bl[20894], bl[20895], bl[20896], bl[20897], bl[20898], bl[20899], bl[20900], bl[20901], bl[20902], bl[20903], bl[20904], bl[20905], bl[20906], bl[20907], bl[20908], bl[20909], bl[20910], bl[20911], bl[20912], bl[20913], bl[20914], bl[20915], bl[20916], bl[20917], bl[20918], bl[20919], bl[20920], bl[20921], bl[20922], bl[20923], bl[20924], bl[20925], bl[20926], bl[20927], bl[20928], bl[20929], bl[20930], bl[20931], bl[20932], bl[20933], bl[20934], bl[20935], bl[20936], bl[20937], bl[20938], bl[20939], bl[20940], bl[20941], bl[20942], bl[20943], bl[20944], bl[20945], bl[20946], bl[20947], bl[20948], bl[20949], bl[20950], bl[20951], bl[20952], bl[20953], bl[20954], bl[20955], bl[20956], bl[20957], bl[20958], bl[20959], bl[20960], bl[20961], bl[20962], bl[20963], bl[20964], bl[20965], bl[20966], bl[20967], bl[20968], bl[20969], bl[20970], bl[20971], bl[20972], bl[20973], bl[20974], bl[20975], bl[20976], bl[20977], bl[20978], bl[20979], bl[20980], bl[20981], bl[20982], bl[20983], bl[20984], bl[20985], bl[20986], bl[20987], bl[20988], bl[20989], bl[20990], bl[20991], bl[20992], bl[20993], bl[20994], bl[20995], bl[20996], bl[20997], bl[20998], bl[20999], bl[21000], bl[21001], bl[21002], bl[21003], bl[21004], bl[21005], bl[21006], bl[21007], bl[21008], bl[21009], bl[21010], bl[21011], bl[21012], bl[21013], bl[21014], bl[21015], bl[21016], bl[21017], bl[21018], bl[21019], bl[21020], bl[21021], bl[21022], bl[21023], bl[21024], bl[21025], bl[21026], bl[21027], bl[21028], bl[21029], bl[21030], bl[21031], bl[21032], bl[21033], bl[21034], bl[21035], bl[21036], bl[21037], bl[21038], bl[21039], bl[21040], bl[21041], bl[21042], bl[21043], bl[21044], bl[21045], bl[21046], bl[21047], bl[21048], bl[21049], bl[21050], bl[21051], bl[21052], bl[21053], bl[21054], bl[21055], bl[21056], bl[21057], bl[21058], bl[21059], bl[21060], bl[21061], bl[21062], bl[21063], bl[21064], bl[21065], bl[21066], bl[21067], bl[21068], bl[21069], bl[21070], bl[21071], bl[21072], bl[21073], bl[21074], bl[21075], bl[21076], bl[21077], bl[21078], bl[21079], bl[21080], bl[21081], bl[21082], bl[21083], bl[21084], bl[21085], bl[21086], bl[21087], bl[21088], bl[21089], bl[21090], bl[21091], bl[21092], bl[21093], bl[21094], bl[21095], bl[21096], bl[21097], bl[21098], bl[21099], bl[21100], bl[21101], bl[21102], bl[21103], bl[21104], bl[21105], bl[21106], bl[21107], bl[21108], bl[21109], bl[21110], bl[21111], bl[21112], bl[21113], bl[21114], bl[21115], bl[21116], bl[21117], bl[21118], bl[21119], bl[21120], bl[21121], bl[21122], bl[21123], bl[21124], bl[21125], bl[21126], bl[21127], bl[21128], bl[21129], bl[21130], bl[21131], bl[21132], bl[21133], bl[21134], bl[21135], bl[21136], bl[21137], bl[21138], bl[21139], bl[21140], bl[21141], bl[21142], bl[21143], bl[21144], bl[21145], bl[21146], bl[21147], bl[21148], bl[21149], bl[21150], bl[21151], bl[21152], bl[21153], bl[21154], bl[21155], bl[21156], bl[21157], bl[21158], bl[21159], bl[21160], bl[21161], bl[21162], bl[21163], bl[21164], bl[21165], bl[21166], bl[21167], bl[21168], bl[21169], bl[21170], bl[21171], bl[21172], bl[21173], bl[21174], bl[21175], bl[21176], bl[21177], bl[21178], bl[21179], bl[21180], bl[21181], bl[21182], bl[21183], bl[21184], bl[21185], bl[21186], bl[21187], bl[21188], bl[21189], bl[21190], bl[21191], bl[21192], bl[21193], bl[21194], bl[21195], bl[21196], bl[21197], bl[21198], bl[21199], bl[21200], bl[21201], bl[21202], bl[21203], bl[21204], bl[21205], bl[21206], bl[21207], bl[21208], bl[21209], bl[21210], bl[21211], bl[21212], bl[21213], bl[21214], bl[21215], bl[21216], bl[21217], bl[21218], bl[21219], bl[21220], bl[21221], bl[21222], bl[21223], bl[21224], bl[21225], bl[21226], bl[21227], bl[21228], bl[21229], bl[21230], bl[21231], bl[21232], bl[21233], bl[21234], bl[21235], bl[21236], bl[21237], bl[21238], bl[21239], bl[21240], bl[21241], bl[21242], bl[21243], bl[21244], bl[21245], bl[21246], bl[21247], bl[21248], bl[21249], bl[21250], bl[21251], bl[21252], bl[21253], bl[21254], bl[21255], bl[21256], bl[21257], bl[21258], bl[21259], bl[21260], bl[21261], bl[21262], bl[21263], bl[21264], bl[21265], bl[21266], bl[21267], bl[21268], bl[21269], bl[21270], bl[21271], bl[21272], bl[21273], bl[21274], bl[21275], bl[21276], bl[21277], bl[21278], bl[21279], bl[21280], bl[21281], bl[21282], bl[21283], bl[21284], bl[21285], bl[21286], bl[21287], bl[21288], bl[21289], bl[21290], bl[21291], bl[21292], bl[21293], bl[21294], bl[21295], bl[21296], bl[21297], bl[21298], bl[21299], bl[21300], bl[21301], bl[21302], bl[21303], bl[21304], bl[21305], bl[21306], bl[21307], bl[21308], bl[21309], bl[21310], bl[21311], bl[21312], bl[21313], bl[21314], bl[21315], bl[21316], bl[21317], bl[21318], bl[21319], bl[21320], bl[21321], bl[21322], bl[21323], bl[21324], bl[21325], bl[21326], bl[21327], bl[21328], bl[21329], bl[21330], bl[21331], bl[21332], bl[21333], bl[21334], bl[21335], bl[21336], bl[21337], bl[21338], bl[21339], bl[21340], bl[21341], bl[21342], bl[21343], bl[21344], bl[21345], bl[21346], bl[21347], bl[21348], bl[21349], bl[21350], bl[21351], bl[21352], bl[21353], bl[21354], bl[21355], bl[21356], bl[21357], bl[21358], bl[21359], bl[21360], bl[21361], bl[21362], bl[21363], bl[21364], bl[21365], bl[21366], bl[21367], bl[21368], bl[21369], bl[21370], bl[21371], bl[21372], bl[21373], bl[21374], bl[21375], bl[21376], bl[21377], bl[21378], bl[21379], bl[21380], bl[21381], bl[21382], bl[21383], bl[21384], bl[21385], bl[21386], bl[21387], bl[21388], bl[21389], bl[21390], bl[21391], bl[21392], bl[21393], bl[21394], bl[21395], bl[21396], bl[21397], bl[21398], bl[21399], bl[21400], bl[21401], bl[21402], bl[21403], bl[21404], bl[21405], bl[21406], bl[21407], bl[21408], bl[21409], bl[21410], bl[21411], bl[21412], bl[21413], bl[21414], bl[21415], bl[21416], bl[21417], bl[21418], bl[21419], bl[21420], bl[21421], bl[21422], bl[21423], bl[21424], bl[21425], bl[21426], bl[21427], bl[21428], bl[21429], bl[21430], bl[21431], bl[21432], bl[21433], bl[21434], bl[21435], bl[21436], bl[21437], bl[21438], bl[21439], bl[21440], bl[21441], bl[21442], bl[21443], bl[21444], bl[21445], bl[21446], bl[21447], bl[21448], bl[21449], bl[21450], bl[21451], bl[21452], bl[21453], bl[21454], bl[21455], bl[21456], bl[21457], bl[21458], bl[21459], bl[21460], bl[21461], bl[21462], bl[21463], bl[21464], bl[21465], bl[21466], bl[21467], bl[21468], bl[21469], bl[21470], bl[21471], bl[21472], bl[21473], bl[21474], bl[21475], bl[21476], bl[21477], bl[21478], bl[21479], bl[21480], bl[21481], bl[21482], bl[21483], bl[21484], bl[21485], bl[21486], bl[21487], bl[21488], bl[21489], bl[21490], bl[21491], bl[21492], bl[21493], bl[21494], bl[21495], bl[21496], bl[21497], bl[21498], bl[21499], bl[21500], bl[21501], bl[21502], bl[21503], bl[21504], bl[21505], bl[21506], bl[21507], bl[696], bl[697], bl[698], bl[699], bl[700], bl[701], bl[702], bl[703], bl[624], bl[625], bl[626], bl[627], bl[628], bl[629], bl[630], bl[631], bl[632], bl[633], bl[634], bl[635], bl[636], bl[637], bl[638], bl[639], bl[640], bl[641], bl[642], bl[643], bl[644], bl[645], bl[646], bl[647], bl[648], bl[649], bl[650], bl[651], bl[652], bl[653], bl[654], bl[655], bl[656], bl[657], bl[658], bl[659], bl[660], bl[661], bl[662], bl[663], bl[664], bl[665], bl[666], bl[667], bl[668], bl[669], bl[670], bl[671], bl[672], bl[673], bl[674], bl[675], bl[676], bl[677], bl[678], bl[679], bl[680], bl[681], bl[682], bl[683], bl[684], bl[685], bl[686], bl[687], bl[688], bl[689], bl[690], bl[691], bl[692], bl[693], bl[694], bl[695], bl[20408], bl[20409], bl[20410], bl[20411], bl[20412], bl[20413], bl[20414], bl[20415], bl[20416], bl[20417], bl[20418], bl[20419], bl[20420], bl[20421], bl[20422], bl[20423], bl[20424], bl[20425], bl[20426], bl[20427], bl[20428], bl[20429], bl[20430], bl[20431], bl[20432], bl[20433], bl[20434], bl[20435], bl[20436], bl[20437], bl[20438], bl[20439], bl[20440], bl[20441], bl[20442], bl[20443], bl[20444], bl[20445], bl[20446], bl[20447], bl[20448], bl[20449], bl[20450], bl[20451], bl[20452], bl[20453], bl[20454], bl[20455], bl[20456], bl[20457], bl[20458], bl[20459], bl[20460], bl[20461], bl[20462], bl[20463], bl[20464], bl[20465], bl[20466], bl[20467], bl[20468], bl[20469], bl[20470], bl[20471], bl[20472], bl[20473], bl[20474], bl[20475], bl[20476], bl[20477], bl[20478], bl[20479], bl[20480], bl[20481], bl[20482], bl[20483], bl[20484], bl[20485], bl[20486], bl[20487], bl[544], bl[545], bl[546], bl[547], bl[548], bl[549], bl[550], bl[551], bl[552], bl[553], bl[554], bl[555], bl[556], bl[557], bl[558], bl[559], bl[560], bl[561], bl[562], bl[563], bl[564], bl[565], bl[566], bl[567], bl[568], bl[569], bl[570], bl[571], bl[572], bl[573], bl[574], bl[575], bl[576], bl[577], bl[578], bl[579], bl[580], bl[581], bl[582], bl[583], bl[584], bl[585], bl[586], bl[587], bl[588], bl[589], bl[590], bl[591], bl[592], bl[593], bl[594], bl[595], bl[596], bl[597], bl[598], bl[599], bl[600], bl[601], bl[602], bl[603], bl[604], bl[605], bl[606], bl[607], bl[608], bl[609], bl[610], bl[611], bl[612], bl[613], bl[614], bl[615], bl[616], bl[617], bl[618], bl[619], bl[620], bl[621], bl[622], bl[623]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    top_tile tile_3__5_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_1__4__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_1__4__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_1__4__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_2__3__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_2__3__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_2__3__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_1__3__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_1__3__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_1__3__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_1__3__grid_top_r_in[1]),
        .grid_left_in(grid_clb_2__4__grid_left_in),
        .grid_bottom_in(grid_clb_2__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[8:15]),
        .io_bottom_in(grid_io_top_2__5__io_bottom_in),
        .chanx_left_in(sb_1__4__0_chanx_right_out),
        .chanx_left_out(cbx_1__4__1_chanx_left_out),
        .chany_bottom_in(sb_1__1__5_chany_top_out),
        .chany_bottom_out(cby_1__1__7_chany_bottom_out),
        .grid_right_out(grid_clb_3__4__grid_left_in),
        .chanx_right_in_0(cbx_1__4__2_chanx_left_out),
        .chanx_right_out_0(sb_1__4__1_chanx_right_out),
        .grid_right_t_inpad(grid_io_top_3__5__io_bottom_in),
        .grid_right_b_in(sb_2__4__grid_right_b_in),
        .grid_bottom_r_in(sb_2__3__grid_top_r_in),
        .grid_bottom_l_in(sb_2__3__grid_top_l_in),
        .grid_left_b_in(sb_1__4__grid_right_b_in),
        .bl({bl[19228], bl[19229], bl[19230], bl[19231], bl[19232], bl[19233], bl[19234], bl[19235], bl[19236], bl[19237], bl[19238], bl[19239], bl[19240], bl[19241], bl[19242], bl[19243], bl[19244], bl[19245], bl[19246], bl[19247], bl[19248], bl[19249], bl[19250], bl[19251], bl[19252], bl[19253], bl[19254], bl[19255], bl[19256], bl[19257], bl[19258], bl[19259], bl[19260], bl[19261], bl[19262], bl[19263], bl[19264], bl[19265], bl[19266], bl[19267], bl[19268], bl[19269], bl[19270], bl[19271], bl[19272], bl[19273], bl[19274], bl[19275], bl[19276], bl[19277], bl[19278], bl[19279], bl[19280], bl[19281], bl[19282], bl[19283], bl[19284], bl[19285], bl[19286], bl[19287], bl[19288], bl[19289], bl[19290], bl[19291], bl[19292], bl[19293], bl[19294], bl[19295], bl[19296], bl[19297], bl[19298], bl[19299], bl[19300], bl[19301], bl[19302], bl[19303], bl[19304], bl[19305], bl[19306], bl[19307], bl[19308], bl[19309], bl[19310], bl[19311], bl[19312], bl[19313], bl[19314], bl[19315], bl[19316], bl[19317], bl[19318], bl[19319], bl[19320], bl[19321], bl[19322], bl[19323], bl[19324], bl[19325], bl[19326], bl[19327], bl[19328], bl[19329], bl[19330], bl[19331], bl[19332], bl[19333], bl[19334], bl[19335], bl[19336], bl[19337], bl[19338], bl[19339], bl[19340], bl[19341], bl[19342], bl[19343], bl[19344], bl[19345], bl[19346], bl[19347], bl[19348], bl[19349], bl[19350], bl[19351], bl[19352], bl[19353], bl[19354], bl[19355], bl[19356], bl[19357], bl[19358], bl[19359], bl[19360], bl[19361], bl[19362], bl[19363], bl[19364], bl[19365], bl[19366], bl[19367], bl[19368], bl[19369], bl[19370], bl[19371], bl[19372], bl[19373], bl[19374], bl[19375], bl[19376], bl[19377], bl[19378], bl[19379], bl[19380], bl[19381], bl[19382], bl[19383], bl[19384], bl[19385], bl[19386], bl[19387], bl[19388], bl[19389], bl[19390], bl[19391], bl[19392], bl[19393], bl[19394], bl[19395], bl[19396], bl[19397], bl[19398], bl[19399], bl[19400], bl[19401], bl[19402], bl[19403], bl[19404], bl[19405], bl[19406], bl[19407], bl[19408], bl[19409], bl[19410], bl[19411], bl[19412], bl[19413], bl[19414], bl[19415], bl[19416], bl[19417], bl[19418], bl[19419], bl[19420], bl[19421], bl[19422], bl[19423], bl[19424], bl[19425], bl[19426], bl[19427], bl[19428], bl[19429], bl[19430], bl[19431], bl[19432], bl[19433], bl[19434], bl[19435], bl[19436], bl[19437], bl[19438], bl[19439], bl[19440], bl[19441], bl[19442], bl[19443], bl[19444], bl[19445], bl[19446], bl[19447], bl[19448], bl[19449], bl[19450], bl[19451], bl[19452], bl[19453], bl[19454], bl[19455], bl[19456], bl[19457], bl[19458], bl[19459], bl[19460], bl[19461], bl[19462], bl[19463], bl[19464], bl[19465], bl[19466], bl[19467], bl[19468], bl[19469], bl[19470], bl[19471], bl[19472], bl[19473], bl[19474], bl[19475], bl[19476], bl[19477], bl[19478], bl[19479], bl[19480], bl[19481], bl[19482], bl[19483], bl[19484], bl[19485], bl[19486], bl[19487], bl[19488], bl[19489], bl[19490], bl[19491], bl[19492], bl[19493], bl[19494], bl[19495], bl[19496], bl[19497], bl[19498], bl[19499], bl[19500], bl[19501], bl[19502], bl[19503], bl[19504], bl[19505], bl[19506], bl[19507], bl[19508], bl[19509], bl[19510], bl[19511], bl[19512], bl[19513], bl[19514], bl[19515], bl[19516], bl[19517], bl[19518], bl[19519], bl[19520], bl[19521], bl[19522], bl[19523], bl[19524], bl[19525], bl[19526], bl[19527], bl[19528], bl[19529], bl[19530], bl[19531], bl[19532], bl[19533], bl[19534], bl[19535], bl[19536], bl[19537], bl[19538], bl[19539], bl[19540], bl[19541], bl[19542], bl[19543], bl[19544], bl[19545], bl[19546], bl[19547], bl[19548], bl[19549], bl[19550], bl[19551], bl[19552], bl[19553], bl[19554], bl[19555], bl[19556], bl[19557], bl[19558], bl[19559], bl[19560], bl[19561], bl[19562], bl[19563], bl[19564], bl[19565], bl[19566], bl[19567], bl[19568], bl[19569], bl[19570], bl[19571], bl[19572], bl[19573], bl[19574], bl[19575], bl[19576], bl[19577], bl[19578], bl[19579], bl[19580], bl[19581], bl[19582], bl[19583], bl[19584], bl[19585], bl[19586], bl[19587], bl[19588], bl[19589], bl[19590], bl[19591], bl[19592], bl[19593], bl[19594], bl[19595], bl[19596], bl[19597], bl[19598], bl[19599], bl[19600], bl[19601], bl[19602], bl[19603], bl[19604], bl[19605], bl[19606], bl[19607], bl[19608], bl[19609], bl[19610], bl[19611], bl[19612], bl[19613], bl[19614], bl[19615], bl[19616], bl[19617], bl[19618], bl[19619], bl[19620], bl[19621], bl[19622], bl[19623], bl[19624], bl[19625], bl[19626], bl[19627], bl[19628], bl[19629], bl[19630], bl[19631], bl[19632], bl[19633], bl[19634], bl[19635], bl[19636], bl[19637], bl[19638], bl[19639], bl[19640], bl[19641], bl[19642], bl[19643], bl[19644], bl[19645], bl[19646], bl[19647], bl[19648], bl[19649], bl[19650], bl[19651], bl[19652], bl[19653], bl[19654], bl[19655], bl[19656], bl[19657], bl[19658], bl[19659], bl[19660], bl[19661], bl[19662], bl[19663], bl[19664], bl[19665], bl[19666], bl[19667], bl[19668], bl[19669], bl[19670], bl[19671], bl[19672], bl[19673], bl[19674], bl[19675], bl[19676], bl[19677], bl[19678], bl[19679], bl[19680], bl[19681], bl[19682], bl[19683], bl[19684], bl[19685], bl[19686], bl[19687], bl[19688], bl[19689], bl[19690], bl[19691], bl[19692], bl[19693], bl[19694], bl[19695], bl[19696], bl[19697], bl[19698], bl[19699], bl[19700], bl[19701], bl[19702], bl[19703], bl[19704], bl[19705], bl[19706], bl[19707], bl[19708], bl[19709], bl[19710], bl[19711], bl[19712], bl[19713], bl[19714], bl[19715], bl[19716], bl[19717], bl[19718], bl[19719], bl[19720], bl[19721], bl[19722], bl[19723], bl[19724], bl[19725], bl[19726], bl[19727], bl[19728], bl[19729], bl[19730], bl[19731], bl[19732], bl[19733], bl[19734], bl[19735], bl[19736], bl[19737], bl[19738], bl[19739], bl[19740], bl[19741], bl[19742], bl[19743], bl[19744], bl[19745], bl[19746], bl[19747], bl[19748], bl[19749], bl[19750], bl[19751], bl[19752], bl[19753], bl[19754], bl[19755], bl[19756], bl[19757], bl[19758], bl[19759], bl[19760], bl[19761], bl[19762], bl[19763], bl[19764], bl[19765], bl[19766], bl[19767], bl[19768], bl[19769], bl[19770], bl[19771], bl[19772], bl[19773], bl[19774], bl[19775], bl[19776], bl[19777], bl[19778], bl[19779], bl[19780], bl[19781], bl[19782], bl[19783], bl[19784], bl[19785], bl[19786], bl[19787], bl[19788], bl[19789], bl[19790], bl[19791], bl[19792], bl[19793], bl[19794], bl[19795], bl[19796], bl[19797], bl[19798], bl[19799], bl[19800], bl[19801], bl[19802], bl[19803], bl[19804], bl[19805], bl[19806], bl[19807], bl[19808], bl[19809], bl[19810], bl[19811], bl[19812], bl[19813], bl[19814], bl[19815], bl[19816], bl[19817], bl[19818], bl[19819], bl[19820], bl[19821], bl[19822], bl[19823], bl[19824], bl[19825], bl[19826], bl[19827], bl[19828], bl[19829], bl[19830], bl[19831], bl[19832], bl[19833], bl[19834], bl[19835], bl[19836], bl[19837], bl[19838], bl[19839], bl[19840], bl[19841], bl[19842], bl[19843], bl[19844], bl[19845], bl[19846], bl[19847], bl[19848], bl[19849], bl[19850], bl[19851], bl[19852], bl[19853], bl[19854], bl[19855], bl[19856], bl[19857], bl[19858], bl[19859], bl[19860], bl[19861], bl[19862], bl[19863], bl[19864], bl[19865], bl[19866], bl[19867], bl[19868], bl[19869], bl[19870], bl[19871], bl[19872], bl[19873], bl[19874], bl[19875], bl[19876], bl[19877], bl[19878], bl[19879], bl[19880], bl[19881], bl[19882], bl[19883], bl[19884], bl[19885], bl[19886], bl[19887], bl[19888], bl[19889], bl[19890], bl[19891], bl[19892], bl[19893], bl[19894], bl[19895], bl[19896], bl[19897], bl[19898], bl[19899], bl[19900], bl[19901], bl[19902], bl[19903], bl[19904], bl[19905], bl[19906], bl[19907], bl[19908], bl[19909], bl[19910], bl[19911], bl[19912], bl[19913], bl[19914], bl[19915], bl[19916], bl[19917], bl[19918], bl[19919], bl[19920], bl[19921], bl[19922], bl[19923], bl[19924], bl[19925], bl[19926], bl[19927], bl[19928], bl[19929], bl[19930], bl[19931], bl[19932], bl[19933], bl[19934], bl[19935], bl[19936], bl[19937], bl[19938], bl[19939], bl[19940], bl[19941], bl[19942], bl[19943], bl[19944], bl[19945], bl[19946], bl[19947], bl[19948], bl[19949], bl[19950], bl[19951], bl[19952], bl[19953], bl[19954], bl[19955], bl[19956], bl[19957], bl[19958], bl[19959], bl[19960], bl[19961], bl[19962], bl[19963], bl[19964], bl[19965], bl[19966], bl[19967], bl[19968], bl[19969], bl[19970], bl[19971], bl[19972], bl[19973], bl[19974], bl[19975], bl[19976], bl[19977], bl[19978], bl[19979], bl[19980], bl[19981], bl[19982], bl[19983], bl[19984], bl[19985], bl[19986], bl[19987], bl[19988], bl[19989], bl[19990], bl[19991], bl[19992], bl[19993], bl[19994], bl[19995], bl[19996], bl[19997], bl[19998], bl[19999], bl[20000], bl[20001], bl[20002], bl[20003], bl[20004], bl[20005], bl[20006], bl[20007], bl[20008], bl[20009], bl[20010], bl[20011], bl[20012], bl[20013], bl[20014], bl[20015], bl[20016], bl[20017], bl[20018], bl[20019], bl[20020], bl[20021], bl[20022], bl[20023], bl[20024], bl[20025], bl[20026], bl[20027], bl[20028], bl[20029], bl[20030], bl[20031], bl[20032], bl[20033], bl[20034], bl[20035], bl[20036], bl[20037], bl[20038], bl[20039], bl[20040], bl[20041], bl[20042], bl[20043], bl[20044], bl[20045], bl[20046], bl[20047], bl[20048], bl[20049], bl[20050], bl[20051], bl[20052], bl[20053], bl[20054], bl[20055], bl[20056], bl[20057], bl[20058], bl[20059], bl[20060], bl[20061], bl[20062], bl[20063], bl[20064], bl[20065], bl[20066], bl[20067], bl[20068], bl[20069], bl[20070], bl[20071], bl[20072], bl[20073], bl[20074], bl[20075], bl[20076], bl[20077], bl[20078], bl[20079], bl[20080], bl[20081], bl[20082], bl[20083], bl[20084], bl[20085], bl[20086], bl[20087], bl[20088], bl[20089], bl[20090], bl[20091], bl[20092], bl[20093], bl[20094], bl[20095], bl[20096], bl[20097], bl[20098], bl[20099], bl[20100], bl[20101], bl[20102], bl[20103], bl[20104], bl[20105], bl[20106], bl[20107], bl[20108], bl[20109], bl[20110], bl[20111], bl[20112], bl[20113], bl[20114], bl[20115], bl[20116], bl[20117], bl[20118], bl[20119], bl[20120], bl[20121], bl[20122], bl[20123], bl[20124], bl[20125], bl[20126], bl[20127], bl[20128], bl[20129], bl[20130], bl[20131], bl[20132], bl[20133], bl[20134], bl[20135], bl[20136], bl[20137], bl[20138], bl[20139], bl[20140], bl[20141], bl[20142], bl[20143], bl[20144], bl[20145], bl[20146], bl[20147], bl[20148], bl[20149], bl[20150], bl[20151], bl[20152], bl[20153], bl[20154], bl[20155], bl[20156], bl[20157], bl[20158], bl[20159], bl[20160], bl[20161], bl[20162], bl[20163], bl[20164], bl[20165], bl[20166], bl[20167], bl[20168], bl[20169], bl[20170], bl[20171], bl[20172], bl[20173], bl[20174], bl[20175], bl[20176], bl[20177], bl[20178], bl[20179], bl[20180], bl[20181], bl[20182], bl[20183], bl[20184], bl[20185], bl[20186], bl[20187], bl[20188], bl[20189], bl[20190], bl[20191], bl[20192], bl[20193], bl[20194], bl[20195], bl[20196], bl[20197], bl[20198], bl[20199], bl[20200], bl[20201], bl[20202], bl[20203], bl[20204], bl[20205], bl[20206], bl[20207], bl[20208], bl[20209], bl[20210], bl[20211], bl[20212], bl[20213], bl[20214], bl[20215], bl[20216], bl[20217], bl[20218], bl[20219], bl[20220], bl[20221], bl[20222], bl[20223], bl[20224], bl[20225], bl[20226], bl[20227], bl[20228], bl[20229], bl[20230], bl[20231], bl[20232], bl[20233], bl[20234], bl[20235], bl[20236], bl[20237], bl[20238], bl[20239], bl[20240], bl[20241], bl[20242], bl[20243], bl[20244], bl[20245], bl[20246], bl[20247], bl[536], bl[537], bl[538], bl[539], bl[540], bl[541], bl[542], bl[543], bl[464], bl[465], bl[466], bl[467], bl[468], bl[469], bl[470], bl[471], bl[472], bl[473], bl[474], bl[475], bl[476], bl[477], bl[478], bl[479], bl[480], bl[481], bl[482], bl[483], bl[484], bl[485], bl[486], bl[487], bl[488], bl[489], bl[490], bl[491], bl[492], bl[493], bl[494], bl[495], bl[496], bl[497], bl[498], bl[499], bl[500], bl[501], bl[502], bl[503], bl[504], bl[505], bl[506], bl[507], bl[508], bl[509], bl[510], bl[511], bl[512], bl[513], bl[514], bl[515], bl[516], bl[517], bl[518], bl[519], bl[520], bl[521], bl[522], bl[523], bl[524], bl[525], bl[526], bl[527], bl[528], bl[529], bl[530], bl[531], bl[532], bl[533], bl[534], bl[535], bl[19148], bl[19149], bl[19150], bl[19151], bl[19152], bl[19153], bl[19154], bl[19155], bl[19156], bl[19157], bl[19158], bl[19159], bl[19160], bl[19161], bl[19162], bl[19163], bl[19164], bl[19165], bl[19166], bl[19167], bl[19168], bl[19169], bl[19170], bl[19171], bl[19172], bl[19173], bl[19174], bl[19175], bl[19176], bl[19177], bl[19178], bl[19179], bl[19180], bl[19181], bl[19182], bl[19183], bl[19184], bl[19185], bl[19186], bl[19187], bl[19188], bl[19189], bl[19190], bl[19191], bl[19192], bl[19193], bl[19194], bl[19195], bl[19196], bl[19197], bl[19198], bl[19199], bl[19200], bl[19201], bl[19202], bl[19203], bl[19204], bl[19205], bl[19206], bl[19207], bl[19208], bl[19209], bl[19210], bl[19211], bl[19212], bl[19213], bl[19214], bl[19215], bl[19216], bl[19217], bl[19218], bl[19219], bl[19220], bl[19221], bl[19222], bl[19223], bl[19224], bl[19225], bl[19226], bl[19227], bl[384], bl[385], bl[386], bl[387], bl[388], bl[389], bl[390], bl[391], bl[392], bl[393], bl[394], bl[395], bl[396], bl[397], bl[398], bl[399], bl[400], bl[401], bl[402], bl[403], bl[404], bl[405], bl[406], bl[407], bl[408], bl[409], bl[410], bl[411], bl[412], bl[413], bl[414], bl[415], bl[416], bl[417], bl[418], bl[419], bl[420], bl[421], bl[422], bl[423], bl[424], bl[425], bl[426], bl[427], bl[428], bl[429], bl[430], bl[431], bl[432], bl[433], bl[434], bl[435], bl[436], bl[437], bl[438], bl[439], bl[440], bl[441], bl[442], bl[443], bl[444], bl[445], bl[446], bl[447], bl[448], bl[449], bl[450], bl[451], bl[452], bl[453], bl[454], bl[455], bl[456], bl[457], bl[458], bl[459], bl[460], bl[461], bl[462], bl[463]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    top_tile tile_4__5_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_2__4__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_2__4__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_2__4__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_3__3__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_3__3__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_3__3__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_2__3__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_2__3__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_2__3__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_2__3__grid_top_r_in[1]),
        .grid_left_in(grid_clb_3__4__grid_left_in),
        .grid_bottom_in(grid_clb_3__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[16:23]),
        .io_bottom_in(grid_io_top_3__5__io_bottom_in),
        .chanx_left_in(sb_1__4__1_chanx_right_out),
        .chanx_left_out(cbx_1__4__2_chanx_left_out),
        .chany_bottom_in(sb_1__1__8_chany_top_out),
        .chany_bottom_out(cby_1__1__11_chany_bottom_out),
        .grid_right_out(grid_clb_4__4__grid_left_in),
        .chanx_right_in_0(cbx_1__4__3_chanx_left_out),
        .chanx_right_out_0(sb_1__4__2_chanx_right_out),
        .grid_right_t_inpad(grid_io_top_4__5__io_bottom_in),
        .grid_right_b_in(sb_3__4__grid_right_b_in),
        .grid_bottom_r_in(sb_3__3__grid_top_r_in),
        .grid_bottom_l_in(sb_3__3__grid_top_l_in),
        .grid_left_b_in(sb_2__4__grid_right_b_in),
        .bl({bl[17968], bl[17969], bl[17970], bl[17971], bl[17972], bl[17973], bl[17974], bl[17975], bl[17976], bl[17977], bl[17978], bl[17979], bl[17980], bl[17981], bl[17982], bl[17983], bl[17984], bl[17985], bl[17986], bl[17987], bl[17988], bl[17989], bl[17990], bl[17991], bl[17992], bl[17993], bl[17994], bl[17995], bl[17996], bl[17997], bl[17998], bl[17999], bl[18000], bl[18001], bl[18002], bl[18003], bl[18004], bl[18005], bl[18006], bl[18007], bl[18008], bl[18009], bl[18010], bl[18011], bl[18012], bl[18013], bl[18014], bl[18015], bl[18016], bl[18017], bl[18018], bl[18019], bl[18020], bl[18021], bl[18022], bl[18023], bl[18024], bl[18025], bl[18026], bl[18027], bl[18028], bl[18029], bl[18030], bl[18031], bl[18032], bl[18033], bl[18034], bl[18035], bl[18036], bl[18037], bl[18038], bl[18039], bl[18040], bl[18041], bl[18042], bl[18043], bl[18044], bl[18045], bl[18046], bl[18047], bl[18048], bl[18049], bl[18050], bl[18051], bl[18052], bl[18053], bl[18054], bl[18055], bl[18056], bl[18057], bl[18058], bl[18059], bl[18060], bl[18061], bl[18062], bl[18063], bl[18064], bl[18065], bl[18066], bl[18067], bl[18068], bl[18069], bl[18070], bl[18071], bl[18072], bl[18073], bl[18074], bl[18075], bl[18076], bl[18077], bl[18078], bl[18079], bl[18080], bl[18081], bl[18082], bl[18083], bl[18084], bl[18085], bl[18086], bl[18087], bl[18088], bl[18089], bl[18090], bl[18091], bl[18092], bl[18093], bl[18094], bl[18095], bl[18096], bl[18097], bl[18098], bl[18099], bl[18100], bl[18101], bl[18102], bl[18103], bl[18104], bl[18105], bl[18106], bl[18107], bl[18108], bl[18109], bl[18110], bl[18111], bl[18112], bl[18113], bl[18114], bl[18115], bl[18116], bl[18117], bl[18118], bl[18119], bl[18120], bl[18121], bl[18122], bl[18123], bl[18124], bl[18125], bl[18126], bl[18127], bl[18128], bl[18129], bl[18130], bl[18131], bl[18132], bl[18133], bl[18134], bl[18135], bl[18136], bl[18137], bl[18138], bl[18139], bl[18140], bl[18141], bl[18142], bl[18143], bl[18144], bl[18145], bl[18146], bl[18147], bl[18148], bl[18149], bl[18150], bl[18151], bl[18152], bl[18153], bl[18154], bl[18155], bl[18156], bl[18157], bl[18158], bl[18159], bl[18160], bl[18161], bl[18162], bl[18163], bl[18164], bl[18165], bl[18166], bl[18167], bl[18168], bl[18169], bl[18170], bl[18171], bl[18172], bl[18173], bl[18174], bl[18175], bl[18176], bl[18177], bl[18178], bl[18179], bl[18180], bl[18181], bl[18182], bl[18183], bl[18184], bl[18185], bl[18186], bl[18187], bl[18188], bl[18189], bl[18190], bl[18191], bl[18192], bl[18193], bl[18194], bl[18195], bl[18196], bl[18197], bl[18198], bl[18199], bl[18200], bl[18201], bl[18202], bl[18203], bl[18204], bl[18205], bl[18206], bl[18207], bl[18208], bl[18209], bl[18210], bl[18211], bl[18212], bl[18213], bl[18214], bl[18215], bl[18216], bl[18217], bl[18218], bl[18219], bl[18220], bl[18221], bl[18222], bl[18223], bl[18224], bl[18225], bl[18226], bl[18227], bl[18228], bl[18229], bl[18230], bl[18231], bl[18232], bl[18233], bl[18234], bl[18235], bl[18236], bl[18237], bl[18238], bl[18239], bl[18240], bl[18241], bl[18242], bl[18243], bl[18244], bl[18245], bl[18246], bl[18247], bl[18248], bl[18249], bl[18250], bl[18251], bl[18252], bl[18253], bl[18254], bl[18255], bl[18256], bl[18257], bl[18258], bl[18259], bl[18260], bl[18261], bl[18262], bl[18263], bl[18264], bl[18265], bl[18266], bl[18267], bl[18268], bl[18269], bl[18270], bl[18271], bl[18272], bl[18273], bl[18274], bl[18275], bl[18276], bl[18277], bl[18278], bl[18279], bl[18280], bl[18281], bl[18282], bl[18283], bl[18284], bl[18285], bl[18286], bl[18287], bl[18288], bl[18289], bl[18290], bl[18291], bl[18292], bl[18293], bl[18294], bl[18295], bl[18296], bl[18297], bl[18298], bl[18299], bl[18300], bl[18301], bl[18302], bl[18303], bl[18304], bl[18305], bl[18306], bl[18307], bl[18308], bl[18309], bl[18310], bl[18311], bl[18312], bl[18313], bl[18314], bl[18315], bl[18316], bl[18317], bl[18318], bl[18319], bl[18320], bl[18321], bl[18322], bl[18323], bl[18324], bl[18325], bl[18326], bl[18327], bl[18328], bl[18329], bl[18330], bl[18331], bl[18332], bl[18333], bl[18334], bl[18335], bl[18336], bl[18337], bl[18338], bl[18339], bl[18340], bl[18341], bl[18342], bl[18343], bl[18344], bl[18345], bl[18346], bl[18347], bl[18348], bl[18349], bl[18350], bl[18351], bl[18352], bl[18353], bl[18354], bl[18355], bl[18356], bl[18357], bl[18358], bl[18359], bl[18360], bl[18361], bl[18362], bl[18363], bl[18364], bl[18365], bl[18366], bl[18367], bl[18368], bl[18369], bl[18370], bl[18371], bl[18372], bl[18373], bl[18374], bl[18375], bl[18376], bl[18377], bl[18378], bl[18379], bl[18380], bl[18381], bl[18382], bl[18383], bl[18384], bl[18385], bl[18386], bl[18387], bl[18388], bl[18389], bl[18390], bl[18391], bl[18392], bl[18393], bl[18394], bl[18395], bl[18396], bl[18397], bl[18398], bl[18399], bl[18400], bl[18401], bl[18402], bl[18403], bl[18404], bl[18405], bl[18406], bl[18407], bl[18408], bl[18409], bl[18410], bl[18411], bl[18412], bl[18413], bl[18414], bl[18415], bl[18416], bl[18417], bl[18418], bl[18419], bl[18420], bl[18421], bl[18422], bl[18423], bl[18424], bl[18425], bl[18426], bl[18427], bl[18428], bl[18429], bl[18430], bl[18431], bl[18432], bl[18433], bl[18434], bl[18435], bl[18436], bl[18437], bl[18438], bl[18439], bl[18440], bl[18441], bl[18442], bl[18443], bl[18444], bl[18445], bl[18446], bl[18447], bl[18448], bl[18449], bl[18450], bl[18451], bl[18452], bl[18453], bl[18454], bl[18455], bl[18456], bl[18457], bl[18458], bl[18459], bl[18460], bl[18461], bl[18462], bl[18463], bl[18464], bl[18465], bl[18466], bl[18467], bl[18468], bl[18469], bl[18470], bl[18471], bl[18472], bl[18473], bl[18474], bl[18475], bl[18476], bl[18477], bl[18478], bl[18479], bl[18480], bl[18481], bl[18482], bl[18483], bl[18484], bl[18485], bl[18486], bl[18487], bl[18488], bl[18489], bl[18490], bl[18491], bl[18492], bl[18493], bl[18494], bl[18495], bl[18496], bl[18497], bl[18498], bl[18499], bl[18500], bl[18501], bl[18502], bl[18503], bl[18504], bl[18505], bl[18506], bl[18507], bl[18508], bl[18509], bl[18510], bl[18511], bl[18512], bl[18513], bl[18514], bl[18515], bl[18516], bl[18517], bl[18518], bl[18519], bl[18520], bl[18521], bl[18522], bl[18523], bl[18524], bl[18525], bl[18526], bl[18527], bl[18528], bl[18529], bl[18530], bl[18531], bl[18532], bl[18533], bl[18534], bl[18535], bl[18536], bl[18537], bl[18538], bl[18539], bl[18540], bl[18541], bl[18542], bl[18543], bl[18544], bl[18545], bl[18546], bl[18547], bl[18548], bl[18549], bl[18550], bl[18551], bl[18552], bl[18553], bl[18554], bl[18555], bl[18556], bl[18557], bl[18558], bl[18559], bl[18560], bl[18561], bl[18562], bl[18563], bl[18564], bl[18565], bl[18566], bl[18567], bl[18568], bl[18569], bl[18570], bl[18571], bl[18572], bl[18573], bl[18574], bl[18575], bl[18576], bl[18577], bl[18578], bl[18579], bl[18580], bl[18581], bl[18582], bl[18583], bl[18584], bl[18585], bl[18586], bl[18587], bl[18588], bl[18589], bl[18590], bl[18591], bl[18592], bl[18593], bl[18594], bl[18595], bl[18596], bl[18597], bl[18598], bl[18599], bl[18600], bl[18601], bl[18602], bl[18603], bl[18604], bl[18605], bl[18606], bl[18607], bl[18608], bl[18609], bl[18610], bl[18611], bl[18612], bl[18613], bl[18614], bl[18615], bl[18616], bl[18617], bl[18618], bl[18619], bl[18620], bl[18621], bl[18622], bl[18623], bl[18624], bl[18625], bl[18626], bl[18627], bl[18628], bl[18629], bl[18630], bl[18631], bl[18632], bl[18633], bl[18634], bl[18635], bl[18636], bl[18637], bl[18638], bl[18639], bl[18640], bl[18641], bl[18642], bl[18643], bl[18644], bl[18645], bl[18646], bl[18647], bl[18648], bl[18649], bl[18650], bl[18651], bl[18652], bl[18653], bl[18654], bl[18655], bl[18656], bl[18657], bl[18658], bl[18659], bl[18660], bl[18661], bl[18662], bl[18663], bl[18664], bl[18665], bl[18666], bl[18667], bl[18668], bl[18669], bl[18670], bl[18671], bl[18672], bl[18673], bl[18674], bl[18675], bl[18676], bl[18677], bl[18678], bl[18679], bl[18680], bl[18681], bl[18682], bl[18683], bl[18684], bl[18685], bl[18686], bl[18687], bl[18688], bl[18689], bl[18690], bl[18691], bl[18692], bl[18693], bl[18694], bl[18695], bl[18696], bl[18697], bl[18698], bl[18699], bl[18700], bl[18701], bl[18702], bl[18703], bl[18704], bl[18705], bl[18706], bl[18707], bl[18708], bl[18709], bl[18710], bl[18711], bl[18712], bl[18713], bl[18714], bl[18715], bl[18716], bl[18717], bl[18718], bl[18719], bl[18720], bl[18721], bl[18722], bl[18723], bl[18724], bl[18725], bl[18726], bl[18727], bl[18728], bl[18729], bl[18730], bl[18731], bl[18732], bl[18733], bl[18734], bl[18735], bl[18736], bl[18737], bl[18738], bl[18739], bl[18740], bl[18741], bl[18742], bl[18743], bl[18744], bl[18745], bl[18746], bl[18747], bl[18748], bl[18749], bl[18750], bl[18751], bl[18752], bl[18753], bl[18754], bl[18755], bl[18756], bl[18757], bl[18758], bl[18759], bl[18760], bl[18761], bl[18762], bl[18763], bl[18764], bl[18765], bl[18766], bl[18767], bl[18768], bl[18769], bl[18770], bl[18771], bl[18772], bl[18773], bl[18774], bl[18775], bl[18776], bl[18777], bl[18778], bl[18779], bl[18780], bl[18781], bl[18782], bl[18783], bl[18784], bl[18785], bl[18786], bl[18787], bl[18788], bl[18789], bl[18790], bl[18791], bl[18792], bl[18793], bl[18794], bl[18795], bl[18796], bl[18797], bl[18798], bl[18799], bl[18800], bl[18801], bl[18802], bl[18803], bl[18804], bl[18805], bl[18806], bl[18807], bl[18808], bl[18809], bl[18810], bl[18811], bl[18812], bl[18813], bl[18814], bl[18815], bl[18816], bl[18817], bl[18818], bl[18819], bl[18820], bl[18821], bl[18822], bl[18823], bl[18824], bl[18825], bl[18826], bl[18827], bl[18828], bl[18829], bl[18830], bl[18831], bl[18832], bl[18833], bl[18834], bl[18835], bl[18836], bl[18837], bl[18838], bl[18839], bl[18840], bl[18841], bl[18842], bl[18843], bl[18844], bl[18845], bl[18846], bl[18847], bl[18848], bl[18849], bl[18850], bl[18851], bl[18852], bl[18853], bl[18854], bl[18855], bl[18856], bl[18857], bl[18858], bl[18859], bl[18860], bl[18861], bl[18862], bl[18863], bl[18864], bl[18865], bl[18866], bl[18867], bl[18868], bl[18869], bl[18870], bl[18871], bl[18872], bl[18873], bl[18874], bl[18875], bl[18876], bl[18877], bl[18878], bl[18879], bl[18880], bl[18881], bl[18882], bl[18883], bl[18884], bl[18885], bl[18886], bl[18887], bl[18888], bl[18889], bl[18890], bl[18891], bl[18892], bl[18893], bl[18894], bl[18895], bl[18896], bl[18897], bl[18898], bl[18899], bl[18900], bl[18901], bl[18902], bl[18903], bl[18904], bl[18905], bl[18906], bl[18907], bl[18908], bl[18909], bl[18910], bl[18911], bl[18912], bl[18913], bl[18914], bl[18915], bl[18916], bl[18917], bl[18918], bl[18919], bl[18920], bl[18921], bl[18922], bl[18923], bl[18924], bl[18925], bl[18926], bl[18927], bl[18928], bl[18929], bl[18930], bl[18931], bl[18932], bl[18933], bl[18934], bl[18935], bl[18936], bl[18937], bl[18938], bl[18939], bl[18940], bl[18941], bl[18942], bl[18943], bl[18944], bl[18945], bl[18946], bl[18947], bl[18948], bl[18949], bl[18950], bl[18951], bl[18952], bl[18953], bl[18954], bl[18955], bl[18956], bl[18957], bl[18958], bl[18959], bl[18960], bl[18961], bl[18962], bl[18963], bl[18964], bl[18965], bl[18966], bl[18967], bl[18968], bl[18969], bl[18970], bl[18971], bl[18972], bl[18973], bl[18974], bl[18975], bl[18976], bl[18977], bl[18978], bl[18979], bl[18980], bl[18981], bl[18982], bl[18983], bl[18984], bl[18985], bl[18986], bl[18987], bl[376], bl[377], bl[378], bl[379], bl[380], bl[381], bl[382], bl[383], bl[304], bl[305], bl[306], bl[307], bl[308], bl[309], bl[310], bl[311], bl[312], bl[313], bl[314], bl[315], bl[316], bl[317], bl[318], bl[319], bl[320], bl[321], bl[322], bl[323], bl[324], bl[325], bl[326], bl[327], bl[328], bl[329], bl[330], bl[331], bl[332], bl[333], bl[334], bl[335], bl[336], bl[337], bl[338], bl[339], bl[340], bl[341], bl[342], bl[343], bl[344], bl[345], bl[346], bl[347], bl[348], bl[349], bl[350], bl[351], bl[352], bl[353], bl[354], bl[355], bl[356], bl[357], bl[358], bl[359], bl[360], bl[361], bl[362], bl[363], bl[364], bl[365], bl[366], bl[367], bl[368], bl[369], bl[370], bl[371], bl[372], bl[373], bl[374], bl[375], bl[17888], bl[17889], bl[17890], bl[17891], bl[17892], bl[17893], bl[17894], bl[17895], bl[17896], bl[17897], bl[17898], bl[17899], bl[17900], bl[17901], bl[17902], bl[17903], bl[17904], bl[17905], bl[17906], bl[17907], bl[17908], bl[17909], bl[17910], bl[17911], bl[17912], bl[17913], bl[17914], bl[17915], bl[17916], bl[17917], bl[17918], bl[17919], bl[17920], bl[17921], bl[17922], bl[17923], bl[17924], bl[17925], bl[17926], bl[17927], bl[17928], bl[17929], bl[17930], bl[17931], bl[17932], bl[17933], bl[17934], bl[17935], bl[17936], bl[17937], bl[17938], bl[17939], bl[17940], bl[17941], bl[17942], bl[17943], bl[17944], bl[17945], bl[17946], bl[17947], bl[17948], bl[17949], bl[17950], bl[17951], bl[17952], bl[17953], bl[17954], bl[17955], bl[17956], bl[17957], bl[17958], bl[17959], bl[17960], bl[17961], bl[17962], bl[17963], bl[17964], bl[17965], bl[17966], bl[17967], bl[224], bl[225], bl[226], bl[227], bl[228], bl[229], bl[230], bl[231], bl[232], bl[233], bl[234], bl[235], bl[236], bl[237], bl[238], bl[239], bl[240], bl[241], bl[242], bl[243], bl[244], bl[245], bl[246], bl[247], bl[248], bl[249], bl[250], bl[251], bl[252], bl[253], bl[254], bl[255], bl[256], bl[257], bl[258], bl[259], bl[260], bl[261], bl[262], bl[263], bl[264], bl[265], bl[266], bl[267], bl[268], bl[269], bl[270], bl[271], bl[272], bl[273], bl[274], bl[275], bl[276], bl[277], bl[278], bl[279], bl[280], bl[281], bl[282], bl[283], bl[284], bl[285], bl[286], bl[287], bl[288], bl[289], bl[290], bl[291], bl[292], bl[293], bl[294], bl[295], bl[296], bl[297], bl[298], bl[299], bl[300], bl[301], bl[302], bl[303]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    top_left_tile tile_1__5_
    (
        .chanx_right_in(cbx_1__4__0_chanx_left_out),
        .chanx_right_out(sb_0__4__0_chanx_right_out),
        .grid_right_t_inpad(grid_io_top_1__5__io_bottom_in),
        .grid_right_b_in(sb_0__4__grid_right_b_in),
        .grid_bottom_r_in(sb_0__3__grid_top_r_in),
        .grid_bottom_l_inpad(grid_io_left_0__4__io_right_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[120:127]),
        .chany_bottom_in_0(sb_0__1__2_chany_top_out),
        .chany_bottom_out_0(cby_0__1__3_chany_bottom_out),
        .grid_right_out(grid_clb_1__4__grid_left_in),
        .bl({bl[704], bl[705], bl[706], bl[707], bl[708], bl[709], bl[710], bl[711], bl[712], bl[713], bl[714], bl[715], bl[716], bl[717], bl[718], bl[719], bl[720], bl[721], bl[722], bl[723], bl[724], bl[725], bl[726], bl[727], bl[728], bl[729], bl[730], bl[731], bl[732], bl[733], bl[734], bl[735], bl[736], bl[737], bl[738], bl[739], bl[740], bl[741], bl[742], bl[743], bl[744], bl[745], bl[746], bl[747], bl[748], bl[749], bl[750], bl[751], bl[752], bl[753], bl[754], bl[755], bl[756], bl[757], bl[758], bl[759], bl[760], bl[761], bl[762], bl[763], bl[764], bl[765], bl[766], bl[767], bl[768], bl[769], bl[770], bl[771], bl[772], bl[773], bl[774], bl[775], bl[776], bl[777], bl[778], bl[779], bl[780], bl[781], bl[782], bl[783], bl[934], bl[935], bl[936], bl[937], bl[938], bl[939], bl[940], bl[941], bl[862], bl[863], bl[864], bl[865], bl[866], bl[867], bl[868], bl[869], bl[870], bl[871], bl[872], bl[873], bl[874], bl[875], bl[876], bl[877], bl[878], bl[879], bl[880], bl[881], bl[882], bl[883], bl[884], bl[885], bl[886], bl[887], bl[888], bl[889], bl[890], bl[891], bl[892], bl[893], bl[894], bl[895], bl[896], bl[897], bl[898], bl[899], bl[900], bl[901], bl[902], bl[903], bl[904], bl[905], bl[906], bl[907], bl[908], bl[909], bl[910], bl[911], bl[912], bl[913], bl[914], bl[915], bl[916], bl[917], bl[918], bl[919], bl[920], bl[921], bl[922], bl[923], bl[924], bl[925], bl[926], bl[927], bl[928], bl[929], bl[930], bl[931], bl[932], bl[933]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    top_right_tile tile_5__5_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_3__4__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_3__4__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_3__4__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_4__3__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_4__3__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_4__3__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_3__3__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_3__3__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_3__3__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_3__3__grid_top_r_in[1]),
        .grid_left_in(grid_clb_4__4__grid_left_in),
        .grid_bottom_in(grid_clb_4__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[24:31]),
        .io_bottom_in(grid_io_top_4__5__io_bottom_in),
        .chanx_left_in(sb_1__4__2_chanx_right_out),
        .chanx_left_out(cbx_1__4__3_chanx_left_out),
        .gfpga_pad_GPIO_PAD_0(gfpga_pad_GPIO_PAD[32:39]),
        .io_left_in(grid_io_right_5__4__io_left_in),
        .chany_bottom_in(sb_4__1__2_chany_top_out),
        .chany_bottom_out(cby_4__1__3_chany_bottom_out),
        .grid_bottom_l_in(sb_4__3__grid_top_l_in),
        .grid_left_b_in(sb_3__4__grid_right_b_in),
        .bl({bl[16708], bl[16709], bl[16710], bl[16711], bl[16712], bl[16713], bl[16714], bl[16715], bl[16716], bl[16717], bl[16718], bl[16719], bl[16720], bl[16721], bl[16722], bl[16723], bl[16724], bl[16725], bl[16726], bl[16727], bl[16728], bl[16729], bl[16730], bl[16731], bl[16732], bl[16733], bl[16734], bl[16735], bl[16736], bl[16737], bl[16738], bl[16739], bl[16740], bl[16741], bl[16742], bl[16743], bl[16744], bl[16745], bl[16746], bl[16747], bl[16748], bl[16749], bl[16750], bl[16751], bl[16752], bl[16753], bl[16754], bl[16755], bl[16756], bl[16757], bl[16758], bl[16759], bl[16760], bl[16761], bl[16762], bl[16763], bl[16764], bl[16765], bl[16766], bl[16767], bl[16768], bl[16769], bl[16770], bl[16771], bl[16772], bl[16773], bl[16774], bl[16775], bl[16776], bl[16777], bl[16778], bl[16779], bl[16780], bl[16781], bl[16782], bl[16783], bl[16784], bl[16785], bl[16786], bl[16787], bl[16788], bl[16789], bl[16790], bl[16791], bl[16792], bl[16793], bl[16794], bl[16795], bl[16796], bl[16797], bl[16798], bl[16799], bl[16800], bl[16801], bl[16802], bl[16803], bl[16804], bl[16805], bl[16806], bl[16807], bl[16808], bl[16809], bl[16810], bl[16811], bl[16812], bl[16813], bl[16814], bl[16815], bl[16816], bl[16817], bl[16818], bl[16819], bl[16820], bl[16821], bl[16822], bl[16823], bl[16824], bl[16825], bl[16826], bl[16827], bl[16828], bl[16829], bl[16830], bl[16831], bl[16832], bl[16833], bl[16834], bl[16835], bl[16836], bl[16837], bl[16838], bl[16839], bl[16840], bl[16841], bl[16842], bl[16843], bl[16844], bl[16845], bl[16846], bl[16847], bl[16848], bl[16849], bl[16850], bl[16851], bl[16852], bl[16853], bl[16854], bl[16855], bl[16856], bl[16857], bl[16858], bl[16859], bl[16860], bl[16861], bl[16862], bl[16863], bl[16864], bl[16865], bl[16866], bl[16867], bl[16868], bl[16869], bl[16870], bl[16871], bl[16872], bl[16873], bl[16874], bl[16875], bl[16876], bl[16877], bl[16878], bl[16879], bl[16880], bl[16881], bl[16882], bl[16883], bl[16884], bl[16885], bl[16886], bl[16887], bl[16888], bl[16889], bl[16890], bl[16891], bl[16892], bl[16893], bl[16894], bl[16895], bl[16896], bl[16897], bl[16898], bl[16899], bl[16900], bl[16901], bl[16902], bl[16903], bl[16904], bl[16905], bl[16906], bl[16907], bl[16908], bl[16909], bl[16910], bl[16911], bl[16912], bl[16913], bl[16914], bl[16915], bl[16916], bl[16917], bl[16918], bl[16919], bl[16920], bl[16921], bl[16922], bl[16923], bl[16924], bl[16925], bl[16926], bl[16927], bl[16928], bl[16929], bl[16930], bl[16931], bl[16932], bl[16933], bl[16934], bl[16935], bl[16936], bl[16937], bl[16938], bl[16939], bl[16940], bl[16941], bl[16942], bl[16943], bl[16944], bl[16945], bl[16946], bl[16947], bl[16948], bl[16949], bl[16950], bl[16951], bl[16952], bl[16953], bl[16954], bl[16955], bl[16956], bl[16957], bl[16958], bl[16959], bl[16960], bl[16961], bl[16962], bl[16963], bl[16964], bl[16965], bl[16966], bl[16967], bl[16968], bl[16969], bl[16970], bl[16971], bl[16972], bl[16973], bl[16974], bl[16975], bl[16976], bl[16977], bl[16978], bl[16979], bl[16980], bl[16981], bl[16982], bl[16983], bl[16984], bl[16985], bl[16986], bl[16987], bl[16988], bl[16989], bl[16990], bl[16991], bl[16992], bl[16993], bl[16994], bl[16995], bl[16996], bl[16997], bl[16998], bl[16999], bl[17000], bl[17001], bl[17002], bl[17003], bl[17004], bl[17005], bl[17006], bl[17007], bl[17008], bl[17009], bl[17010], bl[17011], bl[17012], bl[17013], bl[17014], bl[17015], bl[17016], bl[17017], bl[17018], bl[17019], bl[17020], bl[17021], bl[17022], bl[17023], bl[17024], bl[17025], bl[17026], bl[17027], bl[17028], bl[17029], bl[17030], bl[17031], bl[17032], bl[17033], bl[17034], bl[17035], bl[17036], bl[17037], bl[17038], bl[17039], bl[17040], bl[17041], bl[17042], bl[17043], bl[17044], bl[17045], bl[17046], bl[17047], bl[17048], bl[17049], bl[17050], bl[17051], bl[17052], bl[17053], bl[17054], bl[17055], bl[17056], bl[17057], bl[17058], bl[17059], bl[17060], bl[17061], bl[17062], bl[17063], bl[17064], bl[17065], bl[17066], bl[17067], bl[17068], bl[17069], bl[17070], bl[17071], bl[17072], bl[17073], bl[17074], bl[17075], bl[17076], bl[17077], bl[17078], bl[17079], bl[17080], bl[17081], bl[17082], bl[17083], bl[17084], bl[17085], bl[17086], bl[17087], bl[17088], bl[17089], bl[17090], bl[17091], bl[17092], bl[17093], bl[17094], bl[17095], bl[17096], bl[17097], bl[17098], bl[17099], bl[17100], bl[17101], bl[17102], bl[17103], bl[17104], bl[17105], bl[17106], bl[17107], bl[17108], bl[17109], bl[17110], bl[17111], bl[17112], bl[17113], bl[17114], bl[17115], bl[17116], bl[17117], bl[17118], bl[17119], bl[17120], bl[17121], bl[17122], bl[17123], bl[17124], bl[17125], bl[17126], bl[17127], bl[17128], bl[17129], bl[17130], bl[17131], bl[17132], bl[17133], bl[17134], bl[17135], bl[17136], bl[17137], bl[17138], bl[17139], bl[17140], bl[17141], bl[17142], bl[17143], bl[17144], bl[17145], bl[17146], bl[17147], bl[17148], bl[17149], bl[17150], bl[17151], bl[17152], bl[17153], bl[17154], bl[17155], bl[17156], bl[17157], bl[17158], bl[17159], bl[17160], bl[17161], bl[17162], bl[17163], bl[17164], bl[17165], bl[17166], bl[17167], bl[17168], bl[17169], bl[17170], bl[17171], bl[17172], bl[17173], bl[17174], bl[17175], bl[17176], bl[17177], bl[17178], bl[17179], bl[17180], bl[17181], bl[17182], bl[17183], bl[17184], bl[17185], bl[17186], bl[17187], bl[17188], bl[17189], bl[17190], bl[17191], bl[17192], bl[17193], bl[17194], bl[17195], bl[17196], bl[17197], bl[17198], bl[17199], bl[17200], bl[17201], bl[17202], bl[17203], bl[17204], bl[17205], bl[17206], bl[17207], bl[17208], bl[17209], bl[17210], bl[17211], bl[17212], bl[17213], bl[17214], bl[17215], bl[17216], bl[17217], bl[17218], bl[17219], bl[17220], bl[17221], bl[17222], bl[17223], bl[17224], bl[17225], bl[17226], bl[17227], bl[17228], bl[17229], bl[17230], bl[17231], bl[17232], bl[17233], bl[17234], bl[17235], bl[17236], bl[17237], bl[17238], bl[17239], bl[17240], bl[17241], bl[17242], bl[17243], bl[17244], bl[17245], bl[17246], bl[17247], bl[17248], bl[17249], bl[17250], bl[17251], bl[17252], bl[17253], bl[17254], bl[17255], bl[17256], bl[17257], bl[17258], bl[17259], bl[17260], bl[17261], bl[17262], bl[17263], bl[17264], bl[17265], bl[17266], bl[17267], bl[17268], bl[17269], bl[17270], bl[17271], bl[17272], bl[17273], bl[17274], bl[17275], bl[17276], bl[17277], bl[17278], bl[17279], bl[17280], bl[17281], bl[17282], bl[17283], bl[17284], bl[17285], bl[17286], bl[17287], bl[17288], bl[17289], bl[17290], bl[17291], bl[17292], bl[17293], bl[17294], bl[17295], bl[17296], bl[17297], bl[17298], bl[17299], bl[17300], bl[17301], bl[17302], bl[17303], bl[17304], bl[17305], bl[17306], bl[17307], bl[17308], bl[17309], bl[17310], bl[17311], bl[17312], bl[17313], bl[17314], bl[17315], bl[17316], bl[17317], bl[17318], bl[17319], bl[17320], bl[17321], bl[17322], bl[17323], bl[17324], bl[17325], bl[17326], bl[17327], bl[17328], bl[17329], bl[17330], bl[17331], bl[17332], bl[17333], bl[17334], bl[17335], bl[17336], bl[17337], bl[17338], bl[17339], bl[17340], bl[17341], bl[17342], bl[17343], bl[17344], bl[17345], bl[17346], bl[17347], bl[17348], bl[17349], bl[17350], bl[17351], bl[17352], bl[17353], bl[17354], bl[17355], bl[17356], bl[17357], bl[17358], bl[17359], bl[17360], bl[17361], bl[17362], bl[17363], bl[17364], bl[17365], bl[17366], bl[17367], bl[17368], bl[17369], bl[17370], bl[17371], bl[17372], bl[17373], bl[17374], bl[17375], bl[17376], bl[17377], bl[17378], bl[17379], bl[17380], bl[17381], bl[17382], bl[17383], bl[17384], bl[17385], bl[17386], bl[17387], bl[17388], bl[17389], bl[17390], bl[17391], bl[17392], bl[17393], bl[17394], bl[17395], bl[17396], bl[17397], bl[17398], bl[17399], bl[17400], bl[17401], bl[17402], bl[17403], bl[17404], bl[17405], bl[17406], bl[17407], bl[17408], bl[17409], bl[17410], bl[17411], bl[17412], bl[17413], bl[17414], bl[17415], bl[17416], bl[17417], bl[17418], bl[17419], bl[17420], bl[17421], bl[17422], bl[17423], bl[17424], bl[17425], bl[17426], bl[17427], bl[17428], bl[17429], bl[17430], bl[17431], bl[17432], bl[17433], bl[17434], bl[17435], bl[17436], bl[17437], bl[17438], bl[17439], bl[17440], bl[17441], bl[17442], bl[17443], bl[17444], bl[17445], bl[17446], bl[17447], bl[17448], bl[17449], bl[17450], bl[17451], bl[17452], bl[17453], bl[17454], bl[17455], bl[17456], bl[17457], bl[17458], bl[17459], bl[17460], bl[17461], bl[17462], bl[17463], bl[17464], bl[17465], bl[17466], bl[17467], bl[17468], bl[17469], bl[17470], bl[17471], bl[17472], bl[17473], bl[17474], bl[17475], bl[17476], bl[17477], bl[17478], bl[17479], bl[17480], bl[17481], bl[17482], bl[17483], bl[17484], bl[17485], bl[17486], bl[17487], bl[17488], bl[17489], bl[17490], bl[17491], bl[17492], bl[17493], bl[17494], bl[17495], bl[17496], bl[17497], bl[17498], bl[17499], bl[17500], bl[17501], bl[17502], bl[17503], bl[17504], bl[17505], bl[17506], bl[17507], bl[17508], bl[17509], bl[17510], bl[17511], bl[17512], bl[17513], bl[17514], bl[17515], bl[17516], bl[17517], bl[17518], bl[17519], bl[17520], bl[17521], bl[17522], bl[17523], bl[17524], bl[17525], bl[17526], bl[17527], bl[17528], bl[17529], bl[17530], bl[17531], bl[17532], bl[17533], bl[17534], bl[17535], bl[17536], bl[17537], bl[17538], bl[17539], bl[17540], bl[17541], bl[17542], bl[17543], bl[17544], bl[17545], bl[17546], bl[17547], bl[17548], bl[17549], bl[17550], bl[17551], bl[17552], bl[17553], bl[17554], bl[17555], bl[17556], bl[17557], bl[17558], bl[17559], bl[17560], bl[17561], bl[17562], bl[17563], bl[17564], bl[17565], bl[17566], bl[17567], bl[17568], bl[17569], bl[17570], bl[17571], bl[17572], bl[17573], bl[17574], bl[17575], bl[17576], bl[17577], bl[17578], bl[17579], bl[17580], bl[17581], bl[17582], bl[17583], bl[17584], bl[17585], bl[17586], bl[17587], bl[17588], bl[17589], bl[17590], bl[17591], bl[17592], bl[17593], bl[17594], bl[17595], bl[17596], bl[17597], bl[17598], bl[17599], bl[17600], bl[17601], bl[17602], bl[17603], bl[17604], bl[17605], bl[17606], bl[17607], bl[17608], bl[17609], bl[17610], bl[17611], bl[17612], bl[17613], bl[17614], bl[17615], bl[17616], bl[17617], bl[17618], bl[17619], bl[17620], bl[17621], bl[17622], bl[17623], bl[17624], bl[17625], bl[17626], bl[17627], bl[17628], bl[17629], bl[17630], bl[17631], bl[17632], bl[17633], bl[17634], bl[17635], bl[17636], bl[17637], bl[17638], bl[17639], bl[17640], bl[17641], bl[17642], bl[17643], bl[17644], bl[17645], bl[17646], bl[17647], bl[17648], bl[17649], bl[17650], bl[17651], bl[17652], bl[17653], bl[17654], bl[17655], bl[17656], bl[17657], bl[17658], bl[17659], bl[17660], bl[17661], bl[17662], bl[17663], bl[17664], bl[17665], bl[17666], bl[17667], bl[17668], bl[17669], bl[17670], bl[17671], bl[17672], bl[17673], bl[17674], bl[17675], bl[17676], bl[17677], bl[17678], bl[17679], bl[17680], bl[17681], bl[17682], bl[17683], bl[17684], bl[17685], bl[17686], bl[17687], bl[17688], bl[17689], bl[17690], bl[17691], bl[17692], bl[17693], bl[17694], bl[17695], bl[17696], bl[17697], bl[17698], bl[17699], bl[17700], bl[17701], bl[17702], bl[17703], bl[17704], bl[17705], bl[17706], bl[17707], bl[17708], bl[17709], bl[17710], bl[17711], bl[17712], bl[17713], bl[17714], bl[17715], bl[17716], bl[17717], bl[17718], bl[17719], bl[17720], bl[17721], bl[17722], bl[17723], bl[17724], bl[17725], bl[17726], bl[17727], bl[216], bl[217], bl[218], bl[219], bl[220], bl[221], bl[222], bl[223], bl[144], bl[145], bl[146], bl[147], bl[148], bl[149], bl[150], bl[151], bl[152], bl[153], bl[154], bl[155], bl[156], bl[157], bl[158], bl[159], bl[160], bl[161], bl[162], bl[163], bl[164], bl[165], bl[166], bl[167], bl[168], bl[169], bl[170], bl[171], bl[172], bl[173], bl[174], bl[175], bl[176], bl[177], bl[178], bl[179], bl[180], bl[181], bl[182], bl[183], bl[184], bl[185], bl[186], bl[187], bl[188], bl[189], bl[190], bl[191], bl[192], bl[193], bl[194], bl[195], bl[196], bl[197], bl[198], bl[199], bl[200], bl[201], bl[202], bl[203], bl[204], bl[205], bl[206], bl[207], bl[208], bl[209], bl[210], bl[211], bl[212], bl[213], bl[214], bl[215], bl[56], bl[57], bl[58], bl[59], bl[60], bl[61], bl[62], bl[63], bl[16636], bl[16637], bl[16638], bl[16639], bl[16640], bl[16641], bl[16642], bl[16643], bl[16644], bl[16645], bl[16646], bl[16647], bl[16648], bl[16649], bl[16650], bl[16651], bl[16652], bl[16653], bl[16654], bl[16655], bl[16656], bl[16657], bl[16658], bl[16659], bl[16660], bl[16661], bl[16662], bl[16663], bl[16664], bl[16665], bl[16666], bl[16667], bl[16668], bl[16669], bl[16670], bl[16671], bl[16672], bl[16673], bl[16674], bl[16675], bl[16676], bl[16677], bl[16678], bl[16679], bl[16680], bl[16681], bl[16682], bl[16683], bl[16684], bl[16685], bl[16686], bl[16687], bl[16688], bl[16689], bl[16690], bl[16691], bl[16692], bl[16693], bl[16694], bl[16695], bl[16696], bl[16697], bl[16698], bl[16699], bl[16700], bl[16701], bl[16702], bl[16703], bl[16704], bl[16705], bl[16706], bl[16707], bl[64], bl[65], bl[66], bl[67], bl[68], bl[69], bl[70], bl[71], bl[72], bl[73], bl[74], bl[75], bl[76], bl[77], bl[78], bl[79], bl[80], bl[81], bl[82], bl[83], bl[84], bl[85], bl[86], bl[87], bl[88], bl[89], bl[90], bl[91], bl[92], bl[93], bl[94], bl[95], bl[96], bl[97], bl[98], bl[99], bl[100], bl[101], bl[102], bl[103], bl[104], bl[105], bl[106], bl[107], bl[108], bl[109], bl[110], bl[111], bl[112], bl[113], bl[114], bl[115], bl[116], bl[117], bl[118], bl[119], bl[120], bl[121], bl[122], bl[123], bl[124], bl[125], bl[126], bl[127], bl[128], bl[129], bl[130], bl[131], bl[132], bl[133], bl[134], bl[135], bl[136], bl[137], bl[138], bl[139], bl[140], bl[141], bl[142], bl[143]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    bottom_left_tile tile_1__1_
    (
        .chany_top_in(cby_0__1__0_chany_bottom_out),
        .chanx_right_in(cbx_1__0__0_chanx_left_out),
        .chany_top_out(sb_0__0__0_chany_top_out),
        .chanx_right_out(sb_0__0__0_chanx_right_out),
        .grid_top_r_in(sb_0__0__grid_top_r_in),
        .grid_top_l_inpad(grid_io_left_0__1__io_right_in),
        .grid_right_t_in(sb_0__0__grid_right_t_in),
        .grid_right_b_inpad(grid_io_bottom_1__0__io_top_in),
        .bl(bl[1258:1337]),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    bottom_right_tile tile_5__1_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[64:71]),
        .io_top_in(grid_io_bottom_4__0__io_top_in),
        .chanx_left_in(sb_1__0__2_chanx_right_out),
        .chanx_left_out(cbx_1__0__3_chanx_left_out),
        .grid_top_out(grid_clb_4__1__grid_bottom_in),
        .chany_top_in(cby_4__1__0_chany_bottom_out),
        .chany_top_out(sb_4__0__0_chany_top_out),
        .grid_top_r_inpad(grid_io_right_5__1__io_left_in),
        .grid_top_l_in(sb_4__0__grid_top_l_in),
        .grid_left_t_in(sb_3__0__grid_right_t_in),
        .bl({bl[24], bl[25], bl[26], bl[27], bl[28], bl[29], bl[30], bl[31], bl[5248], bl[5249], bl[5250], bl[5251], bl[5252], bl[5253], bl[5254], bl[5255], bl[5256], bl[5257], bl[5258], bl[5259], bl[5260], bl[5261], bl[5262], bl[5263], bl[5264], bl[5265], bl[5266], bl[5267], bl[5268], bl[5269], bl[5270], bl[5271], bl[5272], bl[5273], bl[5274], bl[5275], bl[5276], bl[5277], bl[5278], bl[5279], bl[5280], bl[5281], bl[5282], bl[5283], bl[5284], bl[5285], bl[5286], bl[5287], bl[5288], bl[5289], bl[5290], bl[5291], bl[5292], bl[5293], bl[5294], bl[5295], bl[5296], bl[5297], bl[5298], bl[5299], bl[5300], bl[5301], bl[5302], bl[5303], bl[5304], bl[5305], bl[5306], bl[5307], bl[5308], bl[5309], bl[5310], bl[5311], bl[5312], bl[5313], bl[5314], bl[5315], bl[5316], bl[5317], bl[5318], bl[5319], bl[5168], bl[5169], bl[5170], bl[5171], bl[5172], bl[5173], bl[5174], bl[5175], bl[5176], bl[5177], bl[5178], bl[5179], bl[5180], bl[5181], bl[5182], bl[5183], bl[5184], bl[5185], bl[5186], bl[5187], bl[5188], bl[5189], bl[5190], bl[5191], bl[5192], bl[5193], bl[5194], bl[5195], bl[5196], bl[5197], bl[5198], bl[5199], bl[5200], bl[5201], bl[5202], bl[5203], bl[5204], bl[5205], bl[5206], bl[5207], bl[5208], bl[5209], bl[5210], bl[5211], bl[5212], bl[5213], bl[5214], bl[5215], bl[5216], bl[5217], bl[5218], bl[5219], bl[5220], bl[5221], bl[5222], bl[5223], bl[5224], bl[5225], bl[5226], bl[5227], bl[5228], bl[5229], bl[5230], bl[5231], bl[5232], bl[5233], bl[5234], bl[5235], bl[5236], bl[5237], bl[5238], bl[5239], bl[5240], bl[5241], bl[5242], bl[5243], bl[5244], bl[5245], bl[5246], bl[5247]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    left_tile tile_1__2_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[96:103]),
        .io_right_in(grid_io_left_0__1__io_right_in),
        .chany_bottom_in(sb_0__0__0_chany_top_out),
        .chany_bottom_out(cby_0__1__0_chany_bottom_out),
        .grid_right_out(grid_clb_1__1__grid_left_in),
        .chany_top_in_0(cby_0__1__1_chany_bottom_out),
        .chanx_right_in(cbx_1__1__0_chanx_left_out),
        .chany_top_out_0(sb_0__1__0_chany_top_out),
        .chanx_right_out(sb_0__1__0_chanx_right_out),
        .grid_top_r_in(sb_0__1__grid_top_r_in),
        .grid_top_l_inpad(grid_io_left_0__2__io_right_in),
        .grid_right_t_in(sb_0__1__grid_right_t_in),
        .grid_right_b_in(sb_0__1__grid_right_b_in),
        .grid_bottom_r_in(sb_0__0__grid_top_r_in),
        .bl({bl[1410], bl[1411], bl[1412], bl[1413], bl[1414], bl[1415], bl[1416], bl[1417], bl[1338], bl[1339], bl[1340], bl[1341], bl[1342], bl[1343], bl[1344], bl[1345], bl[1346], bl[1347], bl[1348], bl[1349], bl[1350], bl[1351], bl[1352], bl[1353], bl[1354], bl[1355], bl[1356], bl[1357], bl[1358], bl[1359], bl[1360], bl[1361], bl[1362], bl[1363], bl[1364], bl[1365], bl[1366], bl[1367], bl[1368], bl[1369], bl[1370], bl[1371], bl[1372], bl[1373], bl[1374], bl[1375], bl[1376], bl[1377], bl[1378], bl[1379], bl[1380], bl[1381], bl[1382], bl[1383], bl[1384], bl[1385], bl[1386], bl[1387], bl[1388], bl[1389], bl[1390], bl[1391], bl[1392], bl[1393], bl[1394], bl[1395], bl[1396], bl[1397], bl[1398], bl[1399], bl[1400], bl[1401], bl[1402], bl[1403], bl[1404], bl[1405], bl[1406], bl[1407], bl[1408], bl[1409], bl[1100], bl[1101], bl[1102], bl[1103], bl[1104], bl[1105], bl[1106], bl[1107], bl[1108], bl[1109], bl[1110], bl[1111], bl[1112], bl[1113], bl[1114], bl[1115], bl[1116], bl[1117], bl[1118], bl[1119], bl[1120], bl[1121], bl[1122], bl[1123], bl[1124], bl[1125], bl[1126], bl[1127], bl[1128], bl[1129], bl[1130], bl[1131], bl[1132], bl[1133], bl[1134], bl[1135], bl[1136], bl[1137], bl[1138], bl[1139], bl[1140], bl[1141], bl[1142], bl[1143], bl[1144], bl[1145], bl[1146], bl[1147], bl[1148], bl[1149], bl[1150], bl[1151], bl[1152], bl[1153], bl[1154], bl[1155], bl[1156], bl[1157], bl[1158], bl[1159], bl[1160], bl[1161], bl[1162], bl[1163], bl[1164], bl[1165], bl[1166], bl[1167], bl[1168], bl[1169], bl[1170], bl[1171], bl[1172], bl[1173], bl[1174], bl[1175], bl[1176], bl[1177]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    left_tile tile_1__3_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[104:111]),
        .io_right_in(grid_io_left_0__2__io_right_in),
        .chany_bottom_in(sb_0__1__0_chany_top_out),
        .chany_bottom_out(cby_0__1__1_chany_bottom_out),
        .grid_right_out(grid_clb_1__2__grid_left_in),
        .chany_top_in_0(cby_0__1__2_chany_bottom_out),
        .chanx_right_in(cbx_1__1__1_chanx_left_out),
        .chany_top_out_0(sb_0__1__1_chany_top_out),
        .chanx_right_out(sb_0__1__1_chanx_right_out),
        .grid_top_r_in(sb_0__2__grid_top_r_in),
        .grid_top_l_inpad(grid_io_left_0__3__io_right_in),
        .grid_right_t_in(sb_0__2__grid_right_t_in),
        .grid_right_b_in(sb_0__2__grid_right_b_in),
        .grid_bottom_r_in(sb_0__1__grid_top_r_in),
        .bl({bl[1250], bl[1251], bl[1252], bl[1253], bl[1254], bl[1255], bl[1256], bl[1257], bl[1178], bl[1179], bl[1180], bl[1181], bl[1182], bl[1183], bl[1184], bl[1185], bl[1186], bl[1187], bl[1188], bl[1189], bl[1190], bl[1191], bl[1192], bl[1193], bl[1194], bl[1195], bl[1196], bl[1197], bl[1198], bl[1199], bl[1200], bl[1201], bl[1202], bl[1203], bl[1204], bl[1205], bl[1206], bl[1207], bl[1208], bl[1209], bl[1210], bl[1211], bl[1212], bl[1213], bl[1214], bl[1215], bl[1216], bl[1217], bl[1218], bl[1219], bl[1220], bl[1221], bl[1222], bl[1223], bl[1224], bl[1225], bl[1226], bl[1227], bl[1228], bl[1229], bl[1230], bl[1231], bl[1232], bl[1233], bl[1234], bl[1235], bl[1236], bl[1237], bl[1238], bl[1239], bl[1240], bl[1241], bl[1242], bl[1243], bl[1244], bl[1245], bl[1246], bl[1247], bl[1248], bl[1249], bl[942], bl[943], bl[944], bl[945], bl[946], bl[947], bl[948], bl[949], bl[950], bl[951], bl[952], bl[953], bl[954], bl[955], bl[956], bl[957], bl[958], bl[959], bl[960], bl[961], bl[962], bl[963], bl[964], bl[965], bl[966], bl[967], bl[968], bl[969], bl[970], bl[971], bl[972], bl[973], bl[974], bl[975], bl[976], bl[977], bl[978], bl[979], bl[980], bl[981], bl[982], bl[983], bl[984], bl[985], bl[986], bl[987], bl[988], bl[989], bl[990], bl[991], bl[992], bl[993], bl[994], bl[995], bl[996], bl[997], bl[998], bl[999], bl[1000], bl[1001], bl[1002], bl[1003], bl[1004], bl[1005], bl[1006], bl[1007], bl[1008], bl[1009], bl[1010], bl[1011], bl[1012], bl[1013], bl[1014], bl[1015], bl[1016], bl[1017], bl[1018], bl[1019]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    left_tile tile_1__4_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[112:119]),
        .io_right_in(grid_io_left_0__3__io_right_in),
        .chany_bottom_in(sb_0__1__1_chany_top_out),
        .chany_bottom_out(cby_0__1__2_chany_bottom_out),
        .grid_right_out(grid_clb_1__3__grid_left_in),
        .chany_top_in_0(cby_0__1__3_chany_bottom_out),
        .chanx_right_in(cbx_1__1__2_chanx_left_out),
        .chany_top_out_0(sb_0__1__2_chany_top_out),
        .chanx_right_out(sb_0__1__2_chanx_right_out),
        .grid_top_r_in(sb_0__3__grid_top_r_in),
        .grid_top_l_inpad(grid_io_left_0__4__io_right_in),
        .grid_right_t_in(sb_0__3__grid_right_t_in),
        .grid_right_b_in(sb_0__3__grid_right_b_in),
        .grid_bottom_r_in(sb_0__2__grid_top_r_in),
        .bl({bl[1092], bl[1093], bl[1094], bl[1095], bl[1096], bl[1097], bl[1098], bl[1099], bl[1020], bl[1021], bl[1022], bl[1023], bl[1024], bl[1025], bl[1026], bl[1027], bl[1028], bl[1029], bl[1030], bl[1031], bl[1032], bl[1033], bl[1034], bl[1035], bl[1036], bl[1037], bl[1038], bl[1039], bl[1040], bl[1041], bl[1042], bl[1043], bl[1044], bl[1045], bl[1046], bl[1047], bl[1048], bl[1049], bl[1050], bl[1051], bl[1052], bl[1053], bl[1054], bl[1055], bl[1056], bl[1057], bl[1058], bl[1059], bl[1060], bl[1061], bl[1062], bl[1063], bl[1064], bl[1065], bl[1066], bl[1067], bl[1068], bl[1069], bl[1070], bl[1071], bl[1072], bl[1073], bl[1074], bl[1075], bl[1076], bl[1077], bl[1078], bl[1079], bl[1080], bl[1081], bl[1082], bl[1083], bl[1084], bl[1085], bl[1086], bl[1087], bl[1088], bl[1089], bl[1090], bl[1091], bl[784], bl[785], bl[786], bl[787], bl[788], bl[789], bl[790], bl[791], bl[792], bl[793], bl[794], bl[795], bl[796], bl[797], bl[798], bl[799], bl[800], bl[801], bl[802], bl[803], bl[804], bl[805], bl[806], bl[807], bl[808], bl[809], bl[810], bl[811], bl[812], bl[813], bl[814], bl[815], bl[816], bl[817], bl[818], bl[819], bl[820], bl[821], bl[822], bl[823], bl[824], bl[825], bl[826], bl[827], bl[828], bl[829], bl[830], bl[831], bl[832], bl[833], bl[834], bl[835], bl[836], bl[837], bl[838], bl[839], bl[840], bl[841], bl[842], bl[843], bl[844], bl[845], bl[846], bl[847], bl[848], bl[849], bl[850], bl[851], bl[852], bl[853], bl[854], bl[855], bl[856], bl[857], bl[858], bl[859], bl[860], bl[861]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    bottom_tile tile_2__1_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[88:95]),
        .io_top_in(grid_io_bottom_1__0__io_top_in),
        .chanx_left_in(sb_0__0__0_chanx_right_out),
        .chanx_left_out(cbx_1__0__0_chanx_left_out),
        .grid_top_out(grid_clb_1__1__grid_bottom_in),
        .chany_top_in(cby_1__1__0_chany_bottom_out),
        .chanx_right_in_0(cbx_1__0__1_chanx_left_out),
        .chany_top_out(sb_1__0__0_chany_top_out),
        .chanx_right_out_0(sb_1__0__0_chanx_right_out),
        .grid_top_r_in(sb_1__0__grid_top_r_in),
        .grid_top_l_in(sb_1__0__grid_top_l_in),
        .grid_right_t_in(sb_1__0__grid_right_t_in),
        .grid_right_b_inpad(grid_io_bottom_2__0__io_top_in),
        .grid_left_t_in(sb_0__0__grid_right_t_in),
        .bl({bl[0], bl[1], bl[2], bl[3], bl[4], bl[5], bl[6], bl[7], bl[1496], bl[1497], bl[1498], bl[1499], bl[1500], bl[1501], bl[1502], bl[1503], bl[1504], bl[1505], bl[1506], bl[1507], bl[1508], bl[1509], bl[1510], bl[1511], bl[1512], bl[1513], bl[1514], bl[1515], bl[1516], bl[1517], bl[1518], bl[1519], bl[1520], bl[1521], bl[1522], bl[1523], bl[1524], bl[1525], bl[1526], bl[1527], bl[1528], bl[1529], bl[1530], bl[1531], bl[1532], bl[1533], bl[1534], bl[1535], bl[1536], bl[1537], bl[1538], bl[1539], bl[1540], bl[1541], bl[1542], bl[1543], bl[1544], bl[1545], bl[1546], bl[1547], bl[1548], bl[1549], bl[1550], bl[1551], bl[1552], bl[1553], bl[1554], bl[1555], bl[1556], bl[1557], bl[1558], bl[1559], bl[1560], bl[1561], bl[1562], bl[1563], bl[1564], bl[1565], bl[1566], bl[1567], bl[1418], bl[1419], bl[1420], bl[1421], bl[1422], bl[1423], bl[1424], bl[1425], bl[1426], bl[1427], bl[1428], bl[1429], bl[1430], bl[1431], bl[1432], bl[1433], bl[1434], bl[1435], bl[1436], bl[1437], bl[1438], bl[1439], bl[1440], bl[1441], bl[1442], bl[1443], bl[1444], bl[1445], bl[1446], bl[1447], bl[1448], bl[1449], bl[1450], bl[1451], bl[1452], bl[1453], bl[1454], bl[1455], bl[1456], bl[1457], bl[1458], bl[1459], bl[1460], bl[1461], bl[1462], bl[1463], bl[1464], bl[1465], bl[1466], bl[1467], bl[1468], bl[1469], bl[1470], bl[1471], bl[1472], bl[1473], bl[1474], bl[1475], bl[1476], bl[1477], bl[1478], bl[1479], bl[1480], bl[1481], bl[1482], bl[1483], bl[1484], bl[1485], bl[1486], bl[1487], bl[1488], bl[1489], bl[1490], bl[1491], bl[1492], bl[1493], bl[1494], bl[1495]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    bottom_tile tile_3__1_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[80:87]),
        .io_top_in(grid_io_bottom_2__0__io_top_in),
        .chanx_left_in(sb_1__0__0_chanx_right_out),
        .chanx_left_out(cbx_1__0__1_chanx_left_out),
        .grid_top_out(grid_clb_2__1__grid_bottom_in),
        .chany_top_in(cby_1__1__4_chany_bottom_out),
        .chanx_right_in_0(cbx_1__0__2_chanx_left_out),
        .chany_top_out(sb_1__0__1_chany_top_out),
        .chanx_right_out_0(sb_1__0__1_chanx_right_out),
        .grid_top_r_in(sb_2__0__grid_top_r_in),
        .grid_top_l_in(sb_2__0__grid_top_l_in),
        .grid_right_t_in(sb_2__0__grid_right_t_in),
        .grid_right_b_inpad(grid_io_bottom_3__0__io_top_in),
        .grid_left_t_in(sb_1__0__grid_right_t_in),
        .bl({bl[8], bl[9], bl[10], bl[11], bl[12], bl[13], bl[14], bl[15], bl[2746], bl[2747], bl[2748], bl[2749], bl[2750], bl[2751], bl[2752], bl[2753], bl[2754], bl[2755], bl[2756], bl[2757], bl[2758], bl[2759], bl[2760], bl[2761], bl[2762], bl[2763], bl[2764], bl[2765], bl[2766], bl[2767], bl[2768], bl[2769], bl[2770], bl[2771], bl[2772], bl[2773], bl[2774], bl[2775], bl[2776], bl[2777], bl[2778], bl[2779], bl[2780], bl[2781], bl[2782], bl[2783], bl[2784], bl[2785], bl[2786], bl[2787], bl[2788], bl[2789], bl[2790], bl[2791], bl[2792], bl[2793], bl[2794], bl[2795], bl[2796], bl[2797], bl[2798], bl[2799], bl[2800], bl[2801], bl[2802], bl[2803], bl[2804], bl[2805], bl[2806], bl[2807], bl[2808], bl[2809], bl[2810], bl[2811], bl[2812], bl[2813], bl[2814], bl[2815], bl[2816], bl[2817], bl[2668], bl[2669], bl[2670], bl[2671], bl[2672], bl[2673], bl[2674], bl[2675], bl[2676], bl[2677], bl[2678], bl[2679], bl[2680], bl[2681], bl[2682], bl[2683], bl[2684], bl[2685], bl[2686], bl[2687], bl[2688], bl[2689], bl[2690], bl[2691], bl[2692], bl[2693], bl[2694], bl[2695], bl[2696], bl[2697], bl[2698], bl[2699], bl[2700], bl[2701], bl[2702], bl[2703], bl[2704], bl[2705], bl[2706], bl[2707], bl[2708], bl[2709], bl[2710], bl[2711], bl[2712], bl[2713], bl[2714], bl[2715], bl[2716], bl[2717], bl[2718], bl[2719], bl[2720], bl[2721], bl[2722], bl[2723], bl[2724], bl[2725], bl[2726], bl[2727], bl[2728], bl[2729], bl[2730], bl[2731], bl[2732], bl[2733], bl[2734], bl[2735], bl[2736], bl[2737], bl[2738], bl[2739], bl[2740], bl[2741], bl[2742], bl[2743], bl[2744], bl[2745]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
    bottom_tile tile_4__1_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[72:79]),
        .io_top_in(grid_io_bottom_3__0__io_top_in),
        .chanx_left_in(sb_1__0__1_chanx_right_out),
        .chanx_left_out(cbx_1__0__2_chanx_left_out),
        .grid_top_out(grid_clb_3__1__grid_bottom_in),
        .chany_top_in(cby_1__1__8_chany_bottom_out),
        .chanx_right_in_0(cbx_1__0__3_chanx_left_out),
        .chany_top_out(sb_1__0__2_chany_top_out),
        .chanx_right_out_0(sb_1__0__2_chanx_right_out),
        .grid_top_r_in(sb_3__0__grid_top_r_in),
        .grid_top_l_in(sb_3__0__grid_top_l_in),
        .grid_right_t_in(sb_3__0__grid_right_t_in),
        .grid_right_b_inpad(grid_io_bottom_4__0__io_top_in),
        .grid_left_t_in(sb_2__0__grid_right_t_in),
        .bl({bl[16], bl[17], bl[18], bl[19], bl[20], bl[21], bl[22], bl[23], bl[3996], bl[3997], bl[3998], bl[3999], bl[4000], bl[4001], bl[4002], bl[4003], bl[4004], bl[4005], bl[4006], bl[4007], bl[4008], bl[4009], bl[4010], bl[4011], bl[4012], bl[4013], bl[4014], bl[4015], bl[4016], bl[4017], bl[4018], bl[4019], bl[4020], bl[4021], bl[4022], bl[4023], bl[4024], bl[4025], bl[4026], bl[4027], bl[4028], bl[4029], bl[4030], bl[4031], bl[4032], bl[4033], bl[4034], bl[4035], bl[4036], bl[4037], bl[4038], bl[4039], bl[4040], bl[4041], bl[4042], bl[4043], bl[4044], bl[4045], bl[4046], bl[4047], bl[4048], bl[4049], bl[4050], bl[4051], bl[4052], bl[4053], bl[4054], bl[4055], bl[4056], bl[4057], bl[4058], bl[4059], bl[4060], bl[4061], bl[4062], bl[4063], bl[4064], bl[4065], bl[4066], bl[4067], bl[3918], bl[3919], bl[3920], bl[3921], bl[3922], bl[3923], bl[3924], bl[3925], bl[3926], bl[3927], bl[3928], bl[3929], bl[3930], bl[3931], bl[3932], bl[3933], bl[3934], bl[3935], bl[3936], bl[3937], bl[3938], bl[3939], bl[3940], bl[3941], bl[3942], bl[3943], bl[3944], bl[3945], bl[3946], bl[3947], bl[3948], bl[3949], bl[3950], bl[3951], bl[3952], bl[3953], bl[3954], bl[3955], bl[3956], bl[3957], bl[3958], bl[3959], bl[3960], bl[3961], bl[3962], bl[3963], bl[3964], bl[3965], bl[3966], bl[3967], bl[3968], bl[3969], bl[3970], bl[3971], bl[3972], bl[3973], bl[3974], bl[3975], bl[3976], bl[3977], bl[3978], bl[3979], bl[3980], bl[3981], bl[3982], bl[3983], bl[3984], bl[3985], bl[3986], bl[3987], bl[3988], bl[3989], bl[3990], bl[3991], bl[3992], bl[3993], bl[3994], bl[3995]}),
        .wl(),
        .wl_in(),
        .wl_out(),
        .bl_in(),
        .bl_out()
    );
endmodule

