//Generated from netlist by SpyDrNet
//netlist name: SDN_VERILOG_NETLIST_logical_tile_io_mode_physical__iopad
module fpga_top
(
    reset,
    clk,
    gfpga_pad_GPIO_PAD
);

    input reset;
    input clk;
    inout [0:127]gfpga_pad_GPIO_PAD;

    wire reset;
    wire clk;
    wire [0:127]gfpga_pad_GPIO_PAD;
    wire [0:19]cbx_1__0__0_chanx_left_out;
    wire [0:19]cbx_1__0__0_chanx_right_out;
    wire [0:19]cbx_1__0__1_chanx_left_out;
    wire [0:19]cbx_1__0__1_chanx_right_out;
    wire [0:19]cbx_1__0__2_chanx_left_out;
    wire [0:19]cbx_1__0__2_chanx_right_out;
    wire [0:19]cbx_1__0__3_chanx_left_out;
    wire [0:19]cbx_1__0__3_chanx_right_out;
    wire [0:19]cbx_1__1__0_chanx_left_out;
    wire [0:19]cbx_1__1__0_chanx_right_out;
    wire [0:19]cbx_1__1__10_chanx_left_out;
    wire [0:19]cbx_1__1__10_chanx_right_out;
    wire [0:19]cbx_1__1__11_chanx_left_out;
    wire [0:19]cbx_1__1__11_chanx_right_out;
    wire [0:19]cbx_1__1__1_chanx_left_out;
    wire [0:19]cbx_1__1__1_chanx_right_out;
    wire [0:19]cbx_1__1__2_chanx_left_out;
    wire [0:19]cbx_1__1__2_chanx_right_out;
    wire [0:19]cbx_1__1__3_chanx_left_out;
    wire [0:19]cbx_1__1__3_chanx_right_out;
    wire [0:19]cbx_1__1__4_chanx_left_out;
    wire [0:19]cbx_1__1__4_chanx_right_out;
    wire [0:19]cbx_1__1__5_chanx_left_out;
    wire [0:19]cbx_1__1__5_chanx_right_out;
    wire [0:19]cbx_1__1__6_chanx_left_out;
    wire [0:19]cbx_1__1__6_chanx_right_out;
    wire [0:19]cbx_1__1__7_chanx_left_out;
    wire [0:19]cbx_1__1__7_chanx_right_out;
    wire [0:19]cbx_1__1__8_chanx_left_out;
    wire [0:19]cbx_1__1__8_chanx_right_out;
    wire [0:19]cbx_1__1__9_chanx_left_out;
    wire [0:19]cbx_1__1__9_chanx_right_out;
    wire [0:19]cbx_1__4__0_chanx_left_out;
    wire [0:19]cbx_1__4__0_chanx_right_out;
    wire [0:19]cbx_1__4__1_chanx_left_out;
    wire [0:19]cbx_1__4__1_chanx_right_out;
    wire [0:19]cbx_1__4__2_chanx_left_out;
    wire [0:19]cbx_1__4__2_chanx_right_out;
    wire [0:19]cbx_1__4__3_chanx_left_out;
    wire [0:19]cbx_1__4__3_chanx_right_out;
    wire [0:19]cby_0__1__0_chany_bottom_out;
    wire [0:19]cby_0__1__0_chany_top_out;
    wire [0:19]cby_0__1__1_chany_bottom_out;
    wire [0:19]cby_0__1__1_chany_top_out;
    wire [0:19]cby_0__1__2_chany_bottom_out;
    wire [0:19]cby_0__1__2_chany_top_out;
    wire [0:19]cby_0__1__3_chany_bottom_out;
    wire [0:19]cby_0__1__3_chany_top_out;
    wire [0:19]cby_1__1__0_chany_bottom_out;
    wire [0:19]cby_1__1__0_chany_top_out;
    wire [0:19]cby_1__1__10_chany_bottom_out;
    wire [0:19]cby_1__1__10_chany_top_out;
    wire [0:19]cby_1__1__11_chany_bottom_out;
    wire [0:19]cby_1__1__11_chany_top_out;
    wire [0:19]cby_1__1__1_chany_bottom_out;
    wire [0:19]cby_1__1__1_chany_top_out;
    wire [0:19]cby_1__1__2_chany_bottom_out;
    wire [0:19]cby_1__1__2_chany_top_out;
    wire [0:19]cby_1__1__3_chany_bottom_out;
    wire [0:19]cby_1__1__3_chany_top_out;
    wire [0:19]cby_1__1__4_chany_bottom_out;
    wire [0:19]cby_1__1__4_chany_top_out;
    wire [0:19]cby_1__1__5_chany_bottom_out;
    wire [0:19]cby_1__1__5_chany_top_out;
    wire [0:19]cby_1__1__6_chany_bottom_out;
    wire [0:19]cby_1__1__6_chany_top_out;
    wire [0:19]cby_1__1__7_chany_bottom_out;
    wire [0:19]cby_1__1__7_chany_top_out;
    wire [0:19]cby_1__1__8_chany_bottom_out;
    wire [0:19]cby_1__1__8_chany_top_out;
    wire [0:19]cby_1__1__9_chany_bottom_out;
    wire [0:19]cby_1__1__9_chany_top_out;
    wire [0:19]cby_4__1__0_chany_bottom_out;
    wire [0:19]cby_4__1__0_chany_top_out;
    wire [0:19]cby_4__1__1_chany_bottom_out;
    wire [0:19]cby_4__1__1_chany_top_out;
    wire [0:19]cby_4__1__2_chany_bottom_out;
    wire [0:19]cby_4__1__2_chany_top_out;
    wire [0:19]cby_4__1__3_chany_bottom_out;
    wire [0:19]cby_4__1__3_chany_top_out;
    wire [0:19]sb_0__0__0_chanx_right_out;
    wire [0:19]sb_0__0__0_chany_top_out;
    wire [0:19]sb_0__1__0_chanx_right_out;
    wire [0:19]sb_0__1__0_chany_bottom_out;
    wire [0:19]sb_0__1__0_chany_top_out;
    wire [0:19]sb_0__1__1_chanx_right_out;
    wire [0:19]sb_0__1__1_chany_bottom_out;
    wire [0:19]sb_0__1__1_chany_top_out;
    wire [0:19]sb_0__1__2_chanx_right_out;
    wire [0:19]sb_0__1__2_chany_bottom_out;
    wire [0:19]sb_0__1__2_chany_top_out;
    wire [0:19]sb_0__4__0_chanx_right_out;
    wire [0:19]sb_0__4__0_chany_bottom_out;
    wire [0:19]sb_1__0__0_chanx_left_out;
    wire [0:19]sb_1__0__0_chanx_right_out;
    wire [0:19]sb_1__0__0_chany_top_out;
    wire [0:19]sb_1__0__1_chanx_left_out;
    wire [0:19]sb_1__0__1_chanx_right_out;
    wire [0:19]sb_1__0__1_chany_top_out;
    wire [0:19]sb_1__0__2_chanx_left_out;
    wire [0:19]sb_1__0__2_chanx_right_out;
    wire [0:19]sb_1__0__2_chany_top_out;
    wire [0:19]sb_1__1__0_chanx_left_out;
    wire [0:19]sb_1__1__0_chanx_right_out;
    wire [0:19]sb_1__1__0_chany_bottom_out;
    wire [0:19]sb_1__1__0_chany_top_out;
    wire [0:19]sb_1__1__1_chanx_left_out;
    wire [0:19]sb_1__1__1_chanx_right_out;
    wire [0:19]sb_1__1__1_chany_bottom_out;
    wire [0:19]sb_1__1__1_chany_top_out;
    wire [0:19]sb_1__1__2_chanx_left_out;
    wire [0:19]sb_1__1__2_chanx_right_out;
    wire [0:19]sb_1__1__2_chany_bottom_out;
    wire [0:19]sb_1__1__2_chany_top_out;
    wire [0:19]sb_1__1__3_chanx_left_out;
    wire [0:19]sb_1__1__3_chanx_right_out;
    wire [0:19]sb_1__1__3_chany_bottom_out;
    wire [0:19]sb_1__1__3_chany_top_out;
    wire [0:19]sb_1__1__4_chanx_left_out;
    wire [0:19]sb_1__1__4_chanx_right_out;
    wire [0:19]sb_1__1__4_chany_bottom_out;
    wire [0:19]sb_1__1__4_chany_top_out;
    wire [0:19]sb_1__1__5_chanx_left_out;
    wire [0:19]sb_1__1__5_chanx_right_out;
    wire [0:19]sb_1__1__5_chany_bottom_out;
    wire [0:19]sb_1__1__5_chany_top_out;
    wire [0:19]sb_1__1__6_chanx_left_out;
    wire [0:19]sb_1__1__6_chanx_right_out;
    wire [0:19]sb_1__1__6_chany_bottom_out;
    wire [0:19]sb_1__1__6_chany_top_out;
    wire [0:19]sb_1__1__7_chanx_left_out;
    wire [0:19]sb_1__1__7_chanx_right_out;
    wire [0:19]sb_1__1__7_chany_bottom_out;
    wire [0:19]sb_1__1__7_chany_top_out;
    wire [0:19]sb_1__1__8_chanx_left_out;
    wire [0:19]sb_1__1__8_chanx_right_out;
    wire [0:19]sb_1__1__8_chany_bottom_out;
    wire [0:19]sb_1__1__8_chany_top_out;
    wire [0:19]sb_1__4__0_chanx_left_out;
    wire [0:19]sb_1__4__0_chanx_right_out;
    wire [0:19]sb_1__4__0_chany_bottom_out;
    wire [0:19]sb_1__4__1_chanx_left_out;
    wire [0:19]sb_1__4__1_chanx_right_out;
    wire [0:19]sb_1__4__1_chany_bottom_out;
    wire [0:19]sb_1__4__2_chanx_left_out;
    wire [0:19]sb_1__4__2_chanx_right_out;
    wire [0:19]sb_1__4__2_chany_bottom_out;
    wire [0:19]sb_4__0__0_chanx_left_out;
    wire [0:19]sb_4__0__0_chany_top_out;
    wire [0:19]sb_4__1__0_chanx_left_out;
    wire [0:19]sb_4__1__0_chany_bottom_out;
    wire [0:19]sb_4__1__0_chany_top_out;
    wire [0:19]sb_4__1__1_chanx_left_out;
    wire [0:19]sb_4__1__1_chany_bottom_out;
    wire [0:19]sb_4__1__1_chany_top_out;
    wire [0:19]sb_4__1__2_chanx_left_out;
    wire [0:19]sb_4__1__2_chany_bottom_out;
    wire [0:19]sb_4__1__2_chany_top_out;
    wire [0:19]sb_4__4__0_chanx_left_out;
    wire [0:19]sb_4__4__0_chany_bottom_out;
    wire [0:9]grid_clb_1__1__grid_left_in;
    wire [0:9]grid_clb_1__1__grid_top_in;
    wire [0:9]grid_clb_1__1__grid_right_in;
    wire [0:9]grid_clb_1__1__grid_bottom_in;
    wire [0:9]grid_clb_1__2__grid_left_in;
    wire [0:9]grid_clb_1__2__grid_top_in;
    wire [0:9]grid_clb_1__2__grid_right_in;
    wire [0:9]grid_clb_1__2__grid_bottom_in;
    wire [0:9]grid_clb_1__3__grid_left_in;
    wire [0:9]grid_clb_1__3__grid_top_in;
    wire [0:9]grid_clb_1__3__grid_right_in;
    wire [0:9]grid_clb_1__3__grid_bottom_in;
    wire [0:9]grid_clb_1__4__grid_left_in;
    wire [0:9]grid_clb_1__4__grid_top_in;
    wire [0:9]grid_clb_1__4__grid_right_in;
    wire [0:9]grid_clb_1__4__grid_bottom_in;
    wire [0:9]grid_clb_2__1__grid_left_in;
    wire [0:9]grid_clb_2__1__grid_top_in;
    wire [0:9]grid_clb_2__1__grid_right_in;
    wire [0:9]grid_clb_2__1__grid_bottom_in;
    wire [0:9]grid_clb_2__2__grid_left_in;
    wire [0:9]grid_clb_2__2__grid_top_in;
    wire [0:9]grid_clb_2__2__grid_right_in;
    wire [0:9]grid_clb_2__2__grid_bottom_in;
    wire [0:9]grid_clb_2__3__grid_left_in;
    wire [0:9]grid_clb_2__3__grid_top_in;
    wire [0:9]grid_clb_2__3__grid_right_in;
    wire [0:9]grid_clb_2__3__grid_bottom_in;
    wire [0:9]grid_clb_2__4__grid_left_in;
    wire [0:9]grid_clb_2__4__grid_top_in;
    wire [0:9]grid_clb_2__4__grid_right_in;
    wire [0:9]grid_clb_2__4__grid_bottom_in;
    wire [0:9]grid_clb_3__1__grid_left_in;
    wire [0:9]grid_clb_3__1__grid_top_in;
    wire [0:9]grid_clb_3__1__grid_right_in;
    wire [0:9]grid_clb_3__1__grid_bottom_in;
    wire [0:9]grid_clb_3__2__grid_left_in;
    wire [0:9]grid_clb_3__2__grid_top_in;
    wire [0:9]grid_clb_3__2__grid_right_in;
    wire [0:9]grid_clb_3__2__grid_bottom_in;
    wire [0:9]grid_clb_3__3__grid_left_in;
    wire [0:9]grid_clb_3__3__grid_top_in;
    wire [0:9]grid_clb_3__3__grid_right_in;
    wire [0:9]grid_clb_3__3__grid_bottom_in;
    wire [0:9]grid_clb_3__4__grid_left_in;
    wire [0:9]grid_clb_3__4__grid_top_in;
    wire [0:9]grid_clb_3__4__grid_right_in;
    wire [0:9]grid_clb_3__4__grid_bottom_in;
    wire [0:9]grid_clb_4__1__grid_left_in;
    wire [0:9]grid_clb_4__1__grid_top_in;
    wire [0:9]grid_clb_4__1__grid_right_in;
    wire [0:9]grid_clb_4__1__grid_bottom_in;
    wire [0:9]grid_clb_4__2__grid_left_in;
    wire [0:9]grid_clb_4__2__grid_top_in;
    wire [0:9]grid_clb_4__2__grid_right_in;
    wire [0:9]grid_clb_4__2__grid_bottom_in;
    wire [0:9]grid_clb_4__3__grid_left_in;
    wire [0:9]grid_clb_4__3__grid_top_in;
    wire [0:9]grid_clb_4__3__grid_right_in;
    wire [0:9]grid_clb_4__3__grid_bottom_in;
    wire [0:9]grid_clb_4__4__grid_left_in;
    wire [0:9]grid_clb_4__4__grid_top_in;
    wire [0:9]grid_clb_4__4__grid_right_in;
    wire [0:9]grid_clb_4__4__grid_bottom_in;
    wire [0:7]grid_io_top_1__5__io_bottom_in;
    wire [0:7]grid_io_top_1__5__io_bottom_out;
    wire [0:7]grid_io_top_2__5__io_bottom_in;
    wire [0:7]grid_io_top_2__5__io_bottom_out;
    wire [0:7]grid_io_top_3__5__io_bottom_in;
    wire [0:7]grid_io_top_3__5__io_bottom_out;
    wire [0:7]grid_io_top_4__5__io_bottom_in;
    wire [0:7]grid_io_top_4__5__io_bottom_out;
    wire [0:7]grid_io_right_5__4__io_left_in;
    wire [0:7]grid_io_right_5__4__io_left_out;
    wire [0:7]grid_io_right_5__3__io_left_in;
    wire [0:7]grid_io_right_5__3__io_left_out;
    wire [0:7]grid_io_right_5__2__io_left_in;
    wire [0:7]grid_io_right_5__2__io_left_out;
    wire [0:7]grid_io_right_5__1__io_left_in;
    wire [0:7]grid_io_right_5__1__io_left_out;
    wire [0:7]grid_io_bottom_4__0__io_top_in;
    wire [0:7]grid_io_bottom_4__0__io_top_out;
    wire [0:7]grid_io_bottom_3__0__io_top_in;
    wire [0:7]grid_io_bottom_3__0__io_top_out;
    wire [0:7]grid_io_bottom_2__0__io_top_in;
    wire [0:7]grid_io_bottom_2__0__io_top_out;
    wire [0:7]grid_io_bottom_1__0__io_top_in;
    wire [0:7]grid_io_bottom_1__0__io_top_out;
    wire [0:7]grid_io_left_0__1__io_right_in;
    wire [0:7]grid_io_left_0__1__io_right_out;
    wire [0:7]grid_io_left_0__2__io_right_in;
    wire [0:7]grid_io_left_0__2__io_right_out;
    wire [0:7]grid_io_left_0__3__io_right_in;
    wire [0:7]grid_io_left_0__3__io_right_out;
    wire [0:7]grid_io_left_0__4__io_right_in;
    wire [0:7]grid_io_left_0__4__io_right_out;
    wire [0:1]sb_0__0__grid_top_r_in;
    wire [0:1]sb_0__0__grid_right_t_in;
    wire [0:1]sb_0__1__grid_top_r_in;
    wire [0:1]sb_0__1__grid_right_t_in;
    wire [0:2]sb_0__1__grid_right_b_in;
    wire [0:1]sb_0__2__grid_top_r_in;
    wire [0:1]sb_0__2__grid_right_t_in;
    wire [0:2]sb_0__2__grid_right_b_in;
    wire [0:1]sb_0__3__grid_top_r_in;
    wire [0:1]sb_0__3__grid_right_t_in;
    wire [0:2]sb_0__3__grid_right_b_in;
    wire [0:2]sb_0__4__grid_right_b_in;
    wire [0:1]sb_1__0__grid_top_r_in;
    wire [0:2]sb_1__0__grid_top_l_in;
    wire [0:1]sb_1__0__grid_right_t_in;
    wire [0:1]sb_2__0__grid_top_r_in;
    wire [0:2]sb_2__0__grid_top_l_in;
    wire [0:1]sb_2__0__grid_right_t_in;
    wire [0:1]sb_3__0__grid_top_r_in;
    wire [0:2]sb_3__0__grid_top_l_in;
    wire [0:1]sb_3__0__grid_right_t_in;
    wire [0:1]sb_1__1__grid_top_r_in;
    wire [0:2]sb_1__1__grid_top_l_in;
    wire [0:1]sb_1__1__grid_right_t_in;
    wire [0:2]sb_1__1__grid_right_b_in;
    wire [0:1]sb_1__2__grid_top_r_in;
    wire [0:2]sb_1__2__grid_top_l_in;
    wire [0:1]sb_1__2__grid_right_t_in;
    wire [0:2]sb_1__2__grid_right_b_in;
    wire [0:1]sb_1__3__grid_top_r_in;
    wire [0:2]sb_1__3__grid_top_l_in;
    wire [0:1]sb_1__3__grid_right_t_in;
    wire [0:2]sb_1__3__grid_right_b_in;
    wire [0:1]sb_2__1__grid_top_r_in;
    wire [0:2]sb_2__1__grid_top_l_in;
    wire [0:1]sb_2__1__grid_right_t_in;
    wire [0:2]sb_2__1__grid_right_b_in;
    wire [0:1]sb_2__2__grid_top_r_in;
    wire [0:2]sb_2__2__grid_top_l_in;
    wire [0:1]sb_2__2__grid_right_t_in;
    wire [0:2]sb_2__2__grid_right_b_in;
    wire [0:1]sb_2__3__grid_top_r_in;
    wire [0:2]sb_2__3__grid_top_l_in;
    wire [0:1]sb_2__3__grid_right_t_in;
    wire [0:2]sb_2__3__grid_right_b_in;
    wire [0:1]sb_3__1__grid_top_r_in;
    wire [0:2]sb_3__1__grid_top_l_in;
    wire [0:1]sb_3__1__grid_right_t_in;
    wire [0:2]sb_3__1__grid_right_b_in;
    wire [0:1]sb_3__2__grid_top_r_in;
    wire [0:2]sb_3__2__grid_top_l_in;
    wire [0:1]sb_3__2__grid_right_t_in;
    wire [0:2]sb_3__2__grid_right_b_in;
    wire [0:1]sb_3__3__grid_top_r_in;
    wire [0:2]sb_3__3__grid_top_l_in;
    wire [0:1]sb_3__3__grid_right_t_in;
    wire [0:2]sb_3__3__grid_right_b_in;
    wire [0:2]sb_1__4__grid_right_b_in;
    wire [0:2]sb_2__4__grid_right_b_in;
    wire [0:2]sb_3__4__grid_right_b_in;
    wire [0:2]sb_4__0__grid_top_l_in;
    wire [0:2]sb_4__1__grid_top_l_in;
    wire [0:2]sb_4__2__grid_top_l_in;
    wire [0:2]sb_4__3__grid_top_l_in;
    wire [19:0]wl_in;
    wire [3:0]tile_1__1__wl_in;
    wire [3:0]tile_2__1__wl_in;
    wire [3:0]tile_3__1__wl_in;
    wire [3:0]tile_4__1__wl_in;
    wire [3:0]tile_5__1__wl_in;
    wire [3:0]tile_1__2__wl_in;
    wire [3:0]tile_2__2__wl_in;
    wire [3:0]tile_3__2__wl_in;
    wire [3:0]tile_4__2__wl_in;
    wire [3:0]tile_5__2__wl_in;
    wire [3:0]tile_1__3__wl_in;
    wire [3:0]tile_2__3__wl_in;
    wire [3:0]tile_3__3__wl_in;
    wire [3:0]tile_4__3__wl_in;
    wire [3:0]tile_5__3__wl_in;
    wire [3:0]tile_1__4__wl_in;
    wire [3:0]tile_2__4__wl_in;
    wire [3:0]tile_3__4__wl_in;
    wire [3:0]tile_4__4__wl_in;
    wire [3:0]tile_5__4__wl_in;
    wire [3:0]tile_1__5__wl_in;
    wire [3:0]tile_2__5__wl_in;
    wire [3:0]tile_3__5__wl_in;
    wire [3:0]tile_4__5__wl_in;
    wire [3:0]tile_5__5__wl_in;
    wire [1299:0]bl_in;
    wire [39:0]tile_1__1__bl_in;
    wire [39:0]tile_1__2__bl_in;
    wire [39:0]tile_1__3__bl_in;
    wire [39:0]tile_1__4__bl_in;
    wire [39:0]tile_1__5__bl_in;
    wire [314:0]tile_2__1__bl_in;
    wire [314:0]tile_2__2__bl_in;
    wire [314:0]tile_2__3__bl_in;
    wire [314:0]tile_2__4__bl_in;
    wire [314:0]tile_2__5__bl_in;
    wire [314:0]tile_3__1__bl_in;
    wire [314:0]tile_3__2__bl_in;
    wire [314:0]tile_3__3__bl_in;
    wire [314:0]tile_3__4__bl_in;
    wire [314:0]tile_3__5__bl_in;
    wire [314:0]tile_4__1__bl_in;
    wire [314:0]tile_4__2__bl_in;
    wire [314:0]tile_4__3__bl_in;
    wire [314:0]tile_4__4__bl_in;
    wire [314:0]tile_4__5__bl_in;
    wire [314:0]tile_5__1__bl_in;
    wire [314:0]tile_5__2__bl_in;
    wire [314:0]tile_5__3__bl_in;
    wire [314:0]tile_5__4__bl_in;
    wire [314:0]tile_5__5__bl_in;

assign tile_1__1__wl_in = wl_in[3:0];
assign tile_1__2__wl_in = wl_in[7:4];
assign tile_1__3__wl_in = wl_in[11:8];
assign tile_1__4__wl_in = wl_in[15:12];
assign tile_1__5__wl_in = wl_in[19:16];
assign tile_1__1__bl_in = bl_in[39:0];
assign tile_2__1__bl_in = bl_in[354:40];
assign tile_3__1__bl_in = bl_in[669:355];
assign tile_4__1__bl_in = bl_in[984:670];
assign tile_5__1__bl_in = bl_in[1299:985];
    tile tile_2__2_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_0__1__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_0__1__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_0__1__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_1__0__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_1__0__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_1__0__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_0__0__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_0__0__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_0__0__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_0__0__grid_top_r_in[1]),
        .grid_left_in(grid_clb_1__1__grid_left_in),
        .grid_bottom_in(grid_clb_1__1__grid_bottom_in),
        .chanx_left_in(sb_0__1__0_chanx_right_out),
        .chanx_left_out(cbx_1__1__0_chanx_left_out),
        .grid_top_out(grid_clb_1__2__grid_bottom_in),
        .chany_bottom_in(sb_1__0__0_chany_top_out),
        .chany_bottom_out(cby_1__1__0_chany_bottom_out),
        .grid_right_out(grid_clb_2__1__grid_left_in),
        .chany_top_in_0(cby_1__1__1_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__3_chanx_left_out),
        .chany_top_out_0(sb_1__1__0_chany_top_out),
        .chanx_right_out_0(sb_1__1__0_chanx_right_out),
        .grid_top_r_in(sb_1__1__grid_top_r_in),
        .grid_top_l_in(sb_1__1__grid_top_l_in),
        .grid_right_t_in(sb_1__1__grid_right_t_in),
        .grid_right_b_in(sb_1__1__grid_right_b_in),
        .grid_bottom_r_in(sb_1__0__grid_top_r_in),
        .grid_bottom_l_in(sb_1__0__grid_top_l_in),
        .grid_left_t_in(sb_0__1__grid_right_t_in),
        .grid_left_b_in(sb_0__1__grid_right_b_in),
        .wl_in(tile_2__2__wl_in),
        .wl_out(tile_3__2__wl_in),
        .bl_in(tile_2__2__bl_in),
        .bl_out(tile_2__3__bl_in)
    );
    tile tile_2__3_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_0__2__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_0__2__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_0__2__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_1__1__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_1__1__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_1__1__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_0__1__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_0__1__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_0__1__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_0__1__grid_top_r_in[1]),
        .grid_left_in(grid_clb_1__2__grid_left_in),
        .grid_bottom_in(grid_clb_1__2__grid_bottom_in),
        .chanx_left_in(sb_0__1__1_chanx_right_out),
        .chanx_left_out(cbx_1__1__1_chanx_left_out),
        .grid_top_out(grid_clb_1__3__grid_bottom_in),
        .chany_bottom_in(sb_1__1__0_chany_top_out),
        .chany_bottom_out(cby_1__1__1_chany_bottom_out),
        .grid_right_out(grid_clb_2__2__grid_left_in),
        .chany_top_in_0(cby_1__1__2_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__4_chanx_left_out),
        .chany_top_out_0(sb_1__1__1_chany_top_out),
        .chanx_right_out_0(sb_1__1__1_chanx_right_out),
        .grid_top_r_in(sb_1__2__grid_top_r_in),
        .grid_top_l_in(sb_1__2__grid_top_l_in),
        .grid_right_t_in(sb_1__2__grid_right_t_in),
        .grid_right_b_in(sb_1__2__grid_right_b_in),
        .grid_bottom_r_in(sb_1__1__grid_top_r_in),
        .grid_bottom_l_in(sb_1__1__grid_top_l_in),
        .grid_left_t_in(sb_0__2__grid_right_t_in),
        .grid_left_b_in(sb_0__2__grid_right_b_in),
        .wl_in(tile_2__3__wl_in),
        .wl_out(tile_3__3__wl_in),
        .bl_in(tile_2__3__bl_in),
        .bl_out(tile_2__4__bl_in)
    );
    tile tile_2__4_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_0__3__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_0__3__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_0__3__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_1__2__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_1__2__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_1__2__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_0__2__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_0__2__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_0__2__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_0__2__grid_top_r_in[1]),
        .grid_left_in(grid_clb_1__3__grid_left_in),
        .grid_bottom_in(grid_clb_1__3__grid_bottom_in),
        .chanx_left_in(sb_0__1__2_chanx_right_out),
        .chanx_left_out(cbx_1__1__2_chanx_left_out),
        .grid_top_out(grid_clb_1__4__grid_bottom_in),
        .chany_bottom_in(sb_1__1__1_chany_top_out),
        .chany_bottom_out(cby_1__1__2_chany_bottom_out),
        .grid_right_out(grid_clb_2__3__grid_left_in),
        .chany_top_in_0(cby_1__1__3_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__5_chanx_left_out),
        .chany_top_out_0(sb_1__1__2_chany_top_out),
        .chanx_right_out_0(sb_1__1__2_chanx_right_out),
        .grid_top_r_in(sb_1__3__grid_top_r_in),
        .grid_top_l_in(sb_1__3__grid_top_l_in),
        .grid_right_t_in(sb_1__3__grid_right_t_in),
        .grid_right_b_in(sb_1__3__grid_right_b_in),
        .grid_bottom_r_in(sb_1__2__grid_top_r_in),
        .grid_bottom_l_in(sb_1__2__grid_top_l_in),
        .grid_left_t_in(sb_0__3__grid_right_t_in),
        .grid_left_b_in(sb_0__3__grid_right_b_in),
        .wl_in(tile_2__4__wl_in),
        .wl_out(tile_3__4__wl_in),
        .bl_in(tile_2__4__bl_in),
        .bl_out(tile_2__5__bl_in)
    );
    tile tile_3__2_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_1__1__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_1__1__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_1__1__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_2__0__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_2__0__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_2__0__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_1__0__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_1__0__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_1__0__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_1__0__grid_top_r_in[1]),
        .grid_left_in(grid_clb_2__1__grid_left_in),
        .grid_bottom_in(grid_clb_2__1__grid_bottom_in),
        .chanx_left_in(sb_1__1__0_chanx_right_out),
        .chanx_left_out(cbx_1__1__3_chanx_left_out),
        .grid_top_out(grid_clb_2__2__grid_bottom_in),
        .chany_bottom_in(sb_1__0__1_chany_top_out),
        .chany_bottom_out(cby_1__1__4_chany_bottom_out),
        .grid_right_out(grid_clb_3__1__grid_left_in),
        .chany_top_in_0(cby_1__1__5_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__6_chanx_left_out),
        .chany_top_out_0(sb_1__1__3_chany_top_out),
        .chanx_right_out_0(sb_1__1__3_chanx_right_out),
        .grid_top_r_in(sb_2__1__grid_top_r_in),
        .grid_top_l_in(sb_2__1__grid_top_l_in),
        .grid_right_t_in(sb_2__1__grid_right_t_in),
        .grid_right_b_in(sb_2__1__grid_right_b_in),
        .grid_bottom_r_in(sb_2__0__grid_top_r_in),
        .grid_bottom_l_in(sb_2__0__grid_top_l_in),
        .grid_left_t_in(sb_1__1__grid_right_t_in),
        .grid_left_b_in(sb_1__1__grid_right_b_in),
        .wl_in(tile_3__2__wl_in),
        .wl_out(tile_4__2__wl_in),
        .bl_in(tile_3__2__bl_in),
        .bl_out(tile_3__3__bl_in)
    );
    tile tile_3__3_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_1__2__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_1__2__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_1__2__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_2__1__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_2__1__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_2__1__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_1__1__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_1__1__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_1__1__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_1__1__grid_top_r_in[1]),
        .grid_left_in(grid_clb_2__2__grid_left_in),
        .grid_bottom_in(grid_clb_2__2__grid_bottom_in),
        .chanx_left_in(sb_1__1__1_chanx_right_out),
        .chanx_left_out(cbx_1__1__4_chanx_left_out),
        .grid_top_out(grid_clb_2__3__grid_bottom_in),
        .chany_bottom_in(sb_1__1__3_chany_top_out),
        .chany_bottom_out(cby_1__1__5_chany_bottom_out),
        .grid_right_out(grid_clb_3__2__grid_left_in),
        .chany_top_in_0(cby_1__1__6_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__7_chanx_left_out),
        .chany_top_out_0(sb_1__1__4_chany_top_out),
        .chanx_right_out_0(sb_1__1__4_chanx_right_out),
        .grid_top_r_in(sb_2__2__grid_top_r_in),
        .grid_top_l_in(sb_2__2__grid_top_l_in),
        .grid_right_t_in(sb_2__2__grid_right_t_in),
        .grid_right_b_in(sb_2__2__grid_right_b_in),
        .grid_bottom_r_in(sb_2__1__grid_top_r_in),
        .grid_bottom_l_in(sb_2__1__grid_top_l_in),
        .grid_left_t_in(sb_1__2__grid_right_t_in),
        .grid_left_b_in(sb_1__2__grid_right_b_in),
        .wl_in(tile_3__3__wl_in),
        .wl_out(tile_4__3__wl_in),
        .bl_in(tile_3__3__bl_in),
        .bl_out(tile_3__4__bl_in)
    );
    tile tile_3__4_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_1__3__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_1__3__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_1__3__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_2__2__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_2__2__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_2__2__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_1__2__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_1__2__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_1__2__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_1__2__grid_top_r_in[1]),
        .grid_left_in(grid_clb_2__3__grid_left_in),
        .grid_bottom_in(grid_clb_2__3__grid_bottom_in),
        .chanx_left_in(sb_1__1__2_chanx_right_out),
        .chanx_left_out(cbx_1__1__5_chanx_left_out),
        .grid_top_out(grid_clb_2__4__grid_bottom_in),
        .chany_bottom_in(sb_1__1__4_chany_top_out),
        .chany_bottom_out(cby_1__1__6_chany_bottom_out),
        .grid_right_out(grid_clb_3__3__grid_left_in),
        .chany_top_in_0(cby_1__1__7_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__8_chanx_left_out),
        .chany_top_out_0(sb_1__1__5_chany_top_out),
        .chanx_right_out_0(sb_1__1__5_chanx_right_out),
        .grid_top_r_in(sb_2__3__grid_top_r_in),
        .grid_top_l_in(sb_2__3__grid_top_l_in),
        .grid_right_t_in(sb_2__3__grid_right_t_in),
        .grid_right_b_in(sb_2__3__grid_right_b_in),
        .grid_bottom_r_in(sb_2__2__grid_top_r_in),
        .grid_bottom_l_in(sb_2__2__grid_top_l_in),
        .grid_left_t_in(sb_1__3__grid_right_t_in),
        .grid_left_b_in(sb_1__3__grid_right_b_in),
        .wl_in(tile_3__4__wl_in),
        .wl_out(tile_4__4__wl_in),
        .bl_in(tile_3__4__bl_in),
        .bl_out(tile_3__5__bl_in)
    );
    tile tile_4__2_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_2__1__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_2__1__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_2__1__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_3__0__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_3__0__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_3__0__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_2__0__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_2__0__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_2__0__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_2__0__grid_top_r_in[1]),
        .grid_left_in(grid_clb_3__1__grid_left_in),
        .grid_bottom_in(grid_clb_3__1__grid_bottom_in),
        .chanx_left_in(sb_1__1__3_chanx_right_out),
        .chanx_left_out(cbx_1__1__6_chanx_left_out),
        .grid_top_out(grid_clb_3__2__grid_bottom_in),
        .chany_bottom_in(sb_1__0__2_chany_top_out),
        .chany_bottom_out(cby_1__1__8_chany_bottom_out),
        .grid_right_out(grid_clb_4__1__grid_left_in),
        .chany_top_in_0(cby_1__1__9_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__9_chanx_left_out),
        .chany_top_out_0(sb_1__1__6_chany_top_out),
        .chanx_right_out_0(sb_1__1__6_chanx_right_out),
        .grid_top_r_in(sb_3__1__grid_top_r_in),
        .grid_top_l_in(sb_3__1__grid_top_l_in),
        .grid_right_t_in(sb_3__1__grid_right_t_in),
        .grid_right_b_in(sb_3__1__grid_right_b_in),
        .grid_bottom_r_in(sb_3__0__grid_top_r_in),
        .grid_bottom_l_in(sb_3__0__grid_top_l_in),
        .grid_left_t_in(sb_2__1__grid_right_t_in),
        .grid_left_b_in(sb_2__1__grid_right_b_in),
        .wl_in(tile_4__2__wl_in),
        .wl_out(tile_5__2__wl_in),
        .bl_in(tile_4__2__bl_in),
        .bl_out(tile_4__3__bl_in)
    );
    tile tile_4__3_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_2__2__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_2__2__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_2__2__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_3__1__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_3__1__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_3__1__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_2__1__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_2__1__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_2__1__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_2__1__grid_top_r_in[1]),
        .grid_left_in(grid_clb_3__2__grid_left_in),
        .grid_bottom_in(grid_clb_3__2__grid_bottom_in),
        .chanx_left_in(sb_1__1__4_chanx_right_out),
        .chanx_left_out(cbx_1__1__7_chanx_left_out),
        .grid_top_out(grid_clb_3__3__grid_bottom_in),
        .chany_bottom_in(sb_1__1__6_chany_top_out),
        .chany_bottom_out(cby_1__1__9_chany_bottom_out),
        .grid_right_out(grid_clb_4__2__grid_left_in),
        .chany_top_in_0(cby_1__1__10_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__10_chanx_left_out),
        .chany_top_out_0(sb_1__1__7_chany_top_out),
        .chanx_right_out_0(sb_1__1__7_chanx_right_out),
        .grid_top_r_in(sb_3__2__grid_top_r_in),
        .grid_top_l_in(sb_3__2__grid_top_l_in),
        .grid_right_t_in(sb_3__2__grid_right_t_in),
        .grid_right_b_in(sb_3__2__grid_right_b_in),
        .grid_bottom_r_in(sb_3__1__grid_top_r_in),
        .grid_bottom_l_in(sb_3__1__grid_top_l_in),
        .grid_left_t_in(sb_2__2__grid_right_t_in),
        .grid_left_b_in(sb_2__2__grid_right_b_in),
        .wl_in(tile_4__3__wl_in),
        .wl_out(tile_5__3__wl_in),
        .bl_in(tile_4__3__bl_in),
        .bl_out(tile_4__4__bl_in)
    );
    tile tile_4__4_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_2__3__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_2__3__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_2__3__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_3__2__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_3__2__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_3__2__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_2__2__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_2__2__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_2__2__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_2__2__grid_top_r_in[1]),
        .grid_left_in(grid_clb_3__3__grid_left_in),
        .grid_bottom_in(grid_clb_3__3__grid_bottom_in),
        .chanx_left_in(sb_1__1__5_chanx_right_out),
        .chanx_left_out(cbx_1__1__8_chanx_left_out),
        .grid_top_out(grid_clb_3__4__grid_bottom_in),
        .chany_bottom_in(sb_1__1__7_chany_top_out),
        .chany_bottom_out(cby_1__1__10_chany_bottom_out),
        .grid_right_out(grid_clb_4__3__grid_left_in),
        .chany_top_in_0(cby_1__1__11_chany_bottom_out),
        .chanx_right_in_0(cbx_1__1__11_chanx_left_out),
        .chany_top_out_0(sb_1__1__8_chany_top_out),
        .chanx_right_out_0(sb_1__1__8_chanx_right_out),
        .grid_top_r_in(sb_3__3__grid_top_r_in),
        .grid_top_l_in(sb_3__3__grid_top_l_in),
        .grid_right_t_in(sb_3__3__grid_right_t_in),
        .grid_right_b_in(sb_3__3__grid_right_b_in),
        .grid_bottom_r_in(sb_3__2__grid_top_r_in),
        .grid_bottom_l_in(sb_3__2__grid_top_l_in),
        .grid_left_t_in(sb_2__3__grid_right_t_in),
        .grid_left_b_in(sb_2__3__grid_right_b_in),
        .wl_in(tile_4__4__wl_in),
        .wl_out(tile_5__4__wl_in),
        .bl_in(tile_4__4__bl_in),
        .bl_out(tile_4__5__bl_in)
    );
    right_tile tile_5__2_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_3__1__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_3__1__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_3__1__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_4__0__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_4__0__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_4__0__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_3__0__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_3__0__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_3__0__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_3__0__grid_top_r_in[1]),
        .grid_left_in(grid_clb_4__1__grid_left_in),
        .grid_bottom_in(grid_clb_4__1__grid_bottom_in),
        .chanx_left_in(sb_1__1__6_chanx_right_out),
        .chanx_left_out(cbx_1__1__9_chanx_left_out),
        .grid_top_out(grid_clb_4__2__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[56:63]),
        .io_left_in(grid_io_right_5__1__io_left_in),
        .chany_bottom_in(sb_4__0__0_chany_top_out),
        .chany_bottom_out(cby_4__1__0_chany_bottom_out),
        .chany_top_in_0(cby_4__1__1_chany_bottom_out),
        .chany_top_out_0(sb_4__1__0_chany_top_out),
        .grid_top_r_inpad(grid_io_right_5__2__io_left_in),
        .grid_top_l_in(sb_4__1__grid_top_l_in),
        .grid_bottom_l_in(sb_4__0__grid_top_l_in),
        .grid_left_t_in(sb_3__1__grid_right_t_in),
        .grid_left_b_in(sb_3__1__grid_right_b_in),
        .wl_in(tile_5__2__wl_in),
        .wl_out(),
        .bl_in(tile_5__2__bl_in),
        .bl_out(tile_5__3__bl_in)
    );
    right_tile tile_5__3_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_3__2__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_3__2__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_3__2__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_4__1__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_4__1__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_4__1__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_3__1__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_3__1__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_3__1__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_3__1__grid_top_r_in[1]),
        .grid_left_in(grid_clb_4__2__grid_left_in),
        .grid_bottom_in(grid_clb_4__2__grid_bottom_in),
        .chanx_left_in(sb_1__1__7_chanx_right_out),
        .chanx_left_out(cbx_1__1__10_chanx_left_out),
        .grid_top_out(grid_clb_4__3__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[48:55]),
        .io_left_in(grid_io_right_5__2__io_left_in),
        .chany_bottom_in(sb_4__1__0_chany_top_out),
        .chany_bottom_out(cby_4__1__1_chany_bottom_out),
        .chany_top_in_0(cby_4__1__2_chany_bottom_out),
        .chany_top_out_0(sb_4__1__1_chany_top_out),
        .grid_top_r_inpad(grid_io_right_5__3__io_left_in),
        .grid_top_l_in(sb_4__2__grid_top_l_in),
        .grid_bottom_l_in(sb_4__1__grid_top_l_in),
        .grid_left_t_in(sb_3__2__grid_right_t_in),
        .grid_left_b_in(sb_3__2__grid_right_b_in),
        .wl_in(tile_5__3__wl_in),
        .wl_out(),
        .bl_in(tile_5__3__bl_in),
        .bl_out(tile_5__4__bl_in)
    );
    right_tile tile_5__4_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_3__3__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_3__3__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_3__3__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_4__2__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_4__2__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_4__2__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_3__2__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_3__2__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_3__2__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_3__2__grid_top_r_in[1]),
        .grid_left_in(grid_clb_4__3__grid_left_in),
        .grid_bottom_in(grid_clb_4__3__grid_bottom_in),
        .chanx_left_in(sb_1__1__8_chanx_right_out),
        .chanx_left_out(cbx_1__1__11_chanx_left_out),
        .grid_top_out(grid_clb_4__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[40:47]),
        .io_left_in(grid_io_right_5__3__io_left_in),
        .chany_bottom_in(sb_4__1__1_chany_top_out),
        .chany_bottom_out(cby_4__1__2_chany_bottom_out),
        .chany_top_in_0(cby_4__1__3_chany_bottom_out),
        .chany_top_out_0(sb_4__1__2_chany_top_out),
        .grid_top_r_inpad(grid_io_right_5__4__io_left_in),
        .grid_top_l_in(sb_4__3__grid_top_l_in),
        .grid_bottom_l_in(sb_4__2__grid_top_l_in),
        .grid_left_t_in(sb_3__3__grid_right_t_in),
        .grid_left_b_in(sb_3__3__grid_right_b_in),
        .wl_in(tile_5__4__wl_in),
        .wl_out(),
        .bl_in(tile_5__4__bl_in),
        .bl_out(tile_5__5__bl_in)
    );
    top_tile tile_2__5_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_0__4__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_0__4__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_0__4__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_1__3__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_1__3__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_1__3__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_0__3__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_0__3__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_0__3__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_0__3__grid_top_r_in[1]),
        .grid_left_in(grid_clb_1__4__grid_left_in),
        .grid_bottom_in(grid_clb_1__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0:7]),
        .io_bottom_in(grid_io_top_1__5__io_bottom_in),
        .chanx_left_in(sb_0__4__0_chanx_right_out),
        .chanx_left_out(cbx_1__4__0_chanx_left_out),
        .chany_bottom_in(sb_1__1__2_chany_top_out),
        .chany_bottom_out(cby_1__1__3_chany_bottom_out),
        .grid_right_out(grid_clb_2__4__grid_left_in),
        .chanx_right_in_0(cbx_1__4__1_chanx_left_out),
        .chanx_right_out_0(sb_1__4__0_chanx_right_out),
        .grid_right_t_inpad(grid_io_top_2__5__io_bottom_in),
        .grid_right_b_in(sb_1__4__grid_right_b_in),
        .grid_bottom_r_in(sb_1__3__grid_top_r_in),
        .grid_bottom_l_in(sb_1__3__grid_top_l_in),
        .grid_left_b_in(sb_0__4__grid_right_b_in),
        .wl_in(tile_2__5__wl_in),
        .wl_out(tile_3__5__wl_in),
        .bl_in(tile_2__5__bl_in),
        .bl_out()
    );
    top_tile tile_3__5_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_1__4__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_1__4__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_1__4__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_2__3__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_2__3__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_2__3__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_1__3__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_1__3__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_1__3__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_1__3__grid_top_r_in[1]),
        .grid_left_in(grid_clb_2__4__grid_left_in),
        .grid_bottom_in(grid_clb_2__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[8:15]),
        .io_bottom_in(grid_io_top_2__5__io_bottom_in),
        .chanx_left_in(sb_1__4__0_chanx_right_out),
        .chanx_left_out(cbx_1__4__1_chanx_left_out),
        .chany_bottom_in(sb_1__1__5_chany_top_out),
        .chany_bottom_out(cby_1__1__7_chany_bottom_out),
        .grid_right_out(grid_clb_3__4__grid_left_in),
        .chanx_right_in_0(cbx_1__4__2_chanx_left_out),
        .chanx_right_out_0(sb_1__4__1_chanx_right_out),
        .grid_right_t_inpad(grid_io_top_3__5__io_bottom_in),
        .grid_right_b_in(sb_2__4__grid_right_b_in),
        .grid_bottom_r_in(sb_2__3__grid_top_r_in),
        .grid_bottom_l_in(sb_2__3__grid_top_l_in),
        .grid_left_b_in(sb_1__4__grid_right_b_in),
        .wl_in(tile_3__5__wl_in),
        .wl_out(tile_4__5__wl_in),
        .bl_in(tile_3__5__bl_in),
        .bl_out()
    );
    top_tile tile_4__5_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_2__4__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_2__4__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_2__4__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_3__3__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_3__3__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_3__3__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_2__3__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_2__3__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_2__3__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_2__3__grid_top_r_in[1]),
        .grid_left_in(grid_clb_3__4__grid_left_in),
        .grid_bottom_in(grid_clb_3__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[16:23]),
        .io_bottom_in(grid_io_top_3__5__io_bottom_in),
        .chanx_left_in(sb_1__4__1_chanx_right_out),
        .chanx_left_out(cbx_1__4__2_chanx_left_out),
        .chany_bottom_in(sb_1__1__8_chany_top_out),
        .chany_bottom_out(cby_1__1__11_chany_bottom_out),
        .grid_right_out(grid_clb_4__4__grid_left_in),
        .chanx_right_in_0(cbx_1__4__3_chanx_left_out),
        .chanx_right_out_0(sb_1__4__2_chanx_right_out),
        .grid_right_t_inpad(grid_io_top_4__5__io_bottom_in),
        .grid_right_b_in(sb_3__4__grid_right_b_in),
        .grid_bottom_r_in(sb_3__3__grid_top_r_in),
        .grid_bottom_l_in(sb_3__3__grid_top_l_in),
        .grid_left_b_in(sb_2__4__grid_right_b_in),
        .wl_in(tile_4__5__wl_in),
        .wl_out(tile_5__5__wl_in),
        .bl_in(tile_4__5__bl_in),
        .bl_out()
    );
    top_left_tile tile_1__5_
    (
        .chanx_right_in(cbx_1__4__0_chanx_left_out),
        .chanx_right_out(sb_0__4__0_chanx_right_out),
        .grid_right_t_inpad(grid_io_top_1__5__io_bottom_in),
        .grid_right_b_in(sb_0__4__grid_right_b_in),
        .grid_bottom_r_in(sb_0__3__grid_top_r_in),
        .grid_bottom_l_inpad(grid_io_left_0__4__io_right_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[120:127]),
        .chany_bottom_in_0(sb_0__1__2_chany_top_out),
        .chany_bottom_out_0(cby_0__1__3_chany_bottom_out),
        .grid_right_out(grid_clb_1__4__grid_left_in),
        .wl_in(tile_1__5__wl_in),
        .wl_out(tile_2__5__wl_in),
        .bl_in(tile_1__5__bl_in),
        .bl_out()
    );
    top_right_tile tile_5__5_
    (
        .reset(reset),
        .clk(clk),
        .bottom_width_0_height_0_subtile_0__pin_clk_0_(),
        .top_width_0_height_0_subtile_0__pin_O_0_(sb_3__4__grid_right_b_in[0]),
        .top_width_0_height_0_subtile_0__pin_O_4_(sb_3__4__grid_right_b_in[1]),
        .top_width_0_height_0_subtile_0__pin_O_8_(sb_3__4__grid_right_b_in[2]),
        .right_width_0_height_0_subtile_0__pin_O_1_(sb_4__3__grid_top_l_in[0]),
        .right_width_0_height_0_subtile_0__pin_O_5_(sb_4__3__grid_top_l_in[1]),
        .right_width_0_height_0_subtile_0__pin_O_9_(sb_4__3__grid_top_l_in[2]),
        .bottom_width_0_height_0_subtile_0__pin_O_2_(sb_3__3__grid_right_t_in[0]),
        .bottom_width_0_height_0_subtile_0__pin_O_6_(sb_3__3__grid_right_t_in[1]),
        .left_width_0_height_0_subtile_0__pin_O_3_(sb_3__3__grid_top_r_in[0]),
        .left_width_0_height_0_subtile_0__pin_O_7_(sb_3__3__grid_top_r_in[1]),
        .grid_left_in(grid_clb_4__4__grid_left_in),
        .grid_bottom_in(grid_clb_4__4__grid_bottom_in),
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[24:31]),
        .io_bottom_in(grid_io_top_4__5__io_bottom_in),
        .chanx_left_in(sb_1__4__2_chanx_right_out),
        .chanx_left_out(cbx_1__4__3_chanx_left_out),
        .gfpga_pad_GPIO_PAD_0(gfpga_pad_GPIO_PAD[32:39]),
        .io_left_in(grid_io_right_5__4__io_left_in),
        .chany_bottom_in(sb_4__1__2_chany_top_out),
        .chany_bottom_out(cby_4__1__3_chany_bottom_out),
        .grid_bottom_l_in(sb_4__3__grid_top_l_in),
        .grid_left_b_in(sb_3__4__grid_right_b_in),
        .wl_in(tile_5__5__wl_in),
        .wl_out(),
        .bl_in(tile_5__5__bl_in),
        .bl_out()
    );
    bottom_left_tile tile_1__1_
    (
        .chany_top_in(cby_0__1__0_chany_bottom_out),
        .chanx_right_in(cbx_1__0__0_chanx_left_out),
        .chany_top_out(sb_0__0__0_chany_top_out),
        .chanx_right_out(sb_0__0__0_chanx_right_out),
        .grid_top_r_in(sb_0__0__grid_top_r_in),
        .grid_top_l_inpad(grid_io_left_0__1__io_right_in),
        .grid_right_t_in(sb_0__0__grid_right_t_in),
        .grid_right_b_inpad(grid_io_bottom_1__0__io_top_in),
        .wl_in(tile_1__1__wl_in),
        .wl_out(tile_2__1__wl_in),
        .bl_in(tile_1__1__bl_in),
        .bl_out(tile_1__2__bl_in)
    );
    bottom_right_tile tile_5__1_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[64:71]),
        .io_top_in(grid_io_bottom_4__0__io_top_in),
        .chanx_left_in(sb_1__0__2_chanx_right_out),
        .chanx_left_out(cbx_1__0__3_chanx_left_out),
        .grid_top_out(grid_clb_4__1__grid_bottom_in),
        .chany_top_in(cby_4__1__0_chany_bottom_out),
        .chany_top_out(sb_4__0__0_chany_top_out),
        .grid_top_r_inpad(grid_io_right_5__1__io_left_in),
        .grid_top_l_in(sb_4__0__grid_top_l_in),
        .grid_left_t_in(sb_3__0__grid_right_t_in),
        .wl_in(tile_5__1__wl_in),
        .wl_out(),
        .bl_in(tile_5__1__bl_in),
        .bl_out(tile_5__2__bl_in)
    );
    left_tile tile_1__2_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[96:103]),
        .io_right_in(grid_io_left_0__1__io_right_in),
        .chany_bottom_in(sb_0__0__0_chany_top_out),
        .chany_bottom_out(cby_0__1__0_chany_bottom_out),
        .grid_right_out(grid_clb_1__1__grid_left_in),
        .chany_top_in_0(cby_0__1__1_chany_bottom_out),
        .chanx_right_in(cbx_1__1__0_chanx_left_out),
        .chany_top_out_0(sb_0__1__0_chany_top_out),
        .chanx_right_out(sb_0__1__0_chanx_right_out),
        .grid_top_r_in(sb_0__1__grid_top_r_in),
        .grid_top_l_inpad(grid_io_left_0__2__io_right_in),
        .grid_right_t_in(sb_0__1__grid_right_t_in),
        .grid_right_b_in(sb_0__1__grid_right_b_in),
        .grid_bottom_r_in(sb_0__0__grid_top_r_in),
        .wl_in(tile_1__2__wl_in),
        .wl_out(tile_2__2__wl_in),
        .bl_in(tile_1__2__bl_in),
        .bl_out(tile_1__3__bl_in)
    );
    left_tile tile_1__3_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[104:111]),
        .io_right_in(grid_io_left_0__2__io_right_in),
        .chany_bottom_in(sb_0__1__0_chany_top_out),
        .chany_bottom_out(cby_0__1__1_chany_bottom_out),
        .grid_right_out(grid_clb_1__2__grid_left_in),
        .chany_top_in_0(cby_0__1__2_chany_bottom_out),
        .chanx_right_in(cbx_1__1__1_chanx_left_out),
        .chany_top_out_0(sb_0__1__1_chany_top_out),
        .chanx_right_out(sb_0__1__1_chanx_right_out),
        .grid_top_r_in(sb_0__2__grid_top_r_in),
        .grid_top_l_inpad(grid_io_left_0__3__io_right_in),
        .grid_right_t_in(sb_0__2__grid_right_t_in),
        .grid_right_b_in(sb_0__2__grid_right_b_in),
        .grid_bottom_r_in(sb_0__1__grid_top_r_in),
        .wl_in(tile_1__3__wl_in),
        .wl_out(tile_2__3__wl_in),
        .bl_in(tile_1__3__bl_in),
        .bl_out(tile_1__4__bl_in)
    );
    left_tile tile_1__4_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[112:119]),
        .io_right_in(grid_io_left_0__3__io_right_in),
        .chany_bottom_in(sb_0__1__1_chany_top_out),
        .chany_bottom_out(cby_0__1__2_chany_bottom_out),
        .grid_right_out(grid_clb_1__3__grid_left_in),
        .chany_top_in_0(cby_0__1__3_chany_bottom_out),
        .chanx_right_in(cbx_1__1__2_chanx_left_out),
        .chany_top_out_0(sb_0__1__2_chany_top_out),
        .chanx_right_out(sb_0__1__2_chanx_right_out),
        .grid_top_r_in(sb_0__3__grid_top_r_in),
        .grid_top_l_inpad(grid_io_left_0__4__io_right_in),
        .grid_right_t_in(sb_0__3__grid_right_t_in),
        .grid_right_b_in(sb_0__3__grid_right_b_in),
        .grid_bottom_r_in(sb_0__2__grid_top_r_in),
        .wl_in(tile_1__4__wl_in),
        .wl_out(tile_2__4__wl_in),
        .bl_in(tile_1__4__bl_in),
        .bl_out(tile_1__5__bl_in)
    );
    bottom_tile tile_2__1_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[88:95]),
        .io_top_in(grid_io_bottom_1__0__io_top_in),
        .chanx_left_in(sb_0__0__0_chanx_right_out),
        .chanx_left_out(cbx_1__0__0_chanx_left_out),
        .grid_top_out(grid_clb_1__1__grid_bottom_in),
        .chany_top_in(cby_1__1__0_chany_bottom_out),
        .chanx_right_in_0(cbx_1__0__1_chanx_left_out),
        .chany_top_out(sb_1__0__0_chany_top_out),
        .chanx_right_out_0(sb_1__0__0_chanx_right_out),
        .grid_top_r_in(sb_1__0__grid_top_r_in),
        .grid_top_l_in(sb_1__0__grid_top_l_in),
        .grid_right_t_in(sb_1__0__grid_right_t_in),
        .grid_right_b_inpad(grid_io_bottom_2__0__io_top_in),
        .grid_left_t_in(sb_0__0__grid_right_t_in),
        .wl_in(tile_2__1__wl_in),
        .wl_out(tile_3__1__wl_in),
        .bl_in(tile_2__1__bl_in),
        .bl_out(tile_2__2__bl_in)
    );
    bottom_tile tile_3__1_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[80:87]),
        .io_top_in(grid_io_bottom_2__0__io_top_in),
        .chanx_left_in(sb_1__0__0_chanx_right_out),
        .chanx_left_out(cbx_1__0__1_chanx_left_out),
        .grid_top_out(grid_clb_2__1__grid_bottom_in),
        .chany_top_in(cby_1__1__4_chany_bottom_out),
        .chanx_right_in_0(cbx_1__0__2_chanx_left_out),
        .chany_top_out(sb_1__0__1_chany_top_out),
        .chanx_right_out_0(sb_1__0__1_chanx_right_out),
        .grid_top_r_in(sb_2__0__grid_top_r_in),
        .grid_top_l_in(sb_2__0__grid_top_l_in),
        .grid_right_t_in(sb_2__0__grid_right_t_in),
        .grid_right_b_inpad(grid_io_bottom_3__0__io_top_in),
        .grid_left_t_in(sb_1__0__grid_right_t_in),
        .wl_in(tile_3__1__wl_in),
        .wl_out(tile_4__1__wl_in),
        .bl_in(tile_3__1__bl_in),
        .bl_out(tile_3__2__bl_in)
    );
    bottom_tile tile_4__1_
    (
        .gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[72:79]),
        .io_top_in(grid_io_bottom_3__0__io_top_in),
        .chanx_left_in(sb_1__0__1_chanx_right_out),
        .chanx_left_out(cbx_1__0__2_chanx_left_out),
        .grid_top_out(grid_clb_3__1__grid_bottom_in),
        .chany_top_in(cby_1__1__8_chany_bottom_out),
        .chanx_right_in_0(cbx_1__0__3_chanx_left_out),
        .chany_top_out(sb_1__0__2_chany_top_out),
        .chanx_right_out_0(sb_1__0__2_chanx_right_out),
        .grid_top_r_in(sb_3__0__grid_top_r_in),
        .grid_top_l_in(sb_3__0__grid_top_l_in),
        .grid_right_t_in(sb_3__0__grid_right_t_in),
        .grid_right_b_inpad(grid_io_bottom_4__0__io_top_in),
        .grid_left_t_in(sb_2__0__grid_right_t_in),
        .wl_in(tile_4__1__wl_in),
        .wl_out(tile_5__1__wl_in),
        .bl_in(tile_4__1__bl_in),
        .bl_out(tile_4__2__bl_in)
    );
endmodule

