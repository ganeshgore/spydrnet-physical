//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Decoders for fabric configuration protocol
//	Organization: University of Utah
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
// `default_nettype wire

// ----- Verilog module for decoder_with_data_in_8to179 -----
module decoder_with_data_in_8to179(enable,
                                   address,
                                   data_in,
                                   data_out);
//----- INPUT PORTS -----
input [0:0] enable;
//----- INPUT PORTS -----
input [0:7] address;
//----- INPUT PORTS -----
input [0:0] data_in;
//----- OUTPUT PORTS -----
output [0:178] data_out;

//----- BEGIN Registered ports -----
reg [0:178] data_out;
//----- END Registered ports -----

// ----- BEGIN Verilog codes for Decoder convert 8-bit addr to 179-bit data -----
always@(address[0:7], enable[0], data_in[0]) begin
	if (enable[0] == 1'b1) begin
		data_out[0:178] = {179{1'bz}};
		case (address[0:7])
			{8{1'b0}} : data_out[0] = data_in[0];
			8'b10000000 : data_out[1] = data_in[0];
			8'b01000000 : data_out[2] = data_in[0];
			8'b11000000 : data_out[3] = data_in[0];
			8'b00100000 : data_out[4] = data_in[0];
			8'b10100000 : data_out[5] = data_in[0];
			8'b01100000 : data_out[6] = data_in[0];
			8'b11100000 : data_out[7] = data_in[0];
			8'b00010000 : data_out[8] = data_in[0];
			8'b10010000 : data_out[9] = data_in[0];
			8'b01010000 : data_out[10] = data_in[0];
			8'b11010000 : data_out[11] = data_in[0];
			8'b00110000 : data_out[12] = data_in[0];
			8'b10110000 : data_out[13] = data_in[0];
			8'b01110000 : data_out[14] = data_in[0];
			8'b11110000 : data_out[15] = data_in[0];
			8'b00001000 : data_out[16] = data_in[0];
			8'b10001000 : data_out[17] = data_in[0];
			8'b01001000 : data_out[18] = data_in[0];
			8'b11001000 : data_out[19] = data_in[0];
			8'b00101000 : data_out[20] = data_in[0];
			8'b10101000 : data_out[21] = data_in[0];
			8'b01101000 : data_out[22] = data_in[0];
			8'b11101000 : data_out[23] = data_in[0];
			8'b00011000 : data_out[24] = data_in[0];
			8'b10011000 : data_out[25] = data_in[0];
			8'b01011000 : data_out[26] = data_in[0];
			8'b11011000 : data_out[27] = data_in[0];
			8'b00111000 : data_out[28] = data_in[0];
			8'b10111000 : data_out[29] = data_in[0];
			8'b01111000 : data_out[30] = data_in[0];
			8'b11111000 : data_out[31] = data_in[0];
			8'b00000100 : data_out[32] = data_in[0];
			8'b10000100 : data_out[33] = data_in[0];
			8'b01000100 : data_out[34] = data_in[0];
			8'b11000100 : data_out[35] = data_in[0];
			8'b00100100 : data_out[36] = data_in[0];
			8'b10100100 : data_out[37] = data_in[0];
			8'b01100100 : data_out[38] = data_in[0];
			8'b11100100 : data_out[39] = data_in[0];
			8'b00010100 : data_out[40] = data_in[0];
			8'b10010100 : data_out[41] = data_in[0];
			8'b01010100 : data_out[42] = data_in[0];
			8'b11010100 : data_out[43] = data_in[0];
			8'b00110100 : data_out[44] = data_in[0];
			8'b10110100 : data_out[45] = data_in[0];
			8'b01110100 : data_out[46] = data_in[0];
			8'b11110100 : data_out[47] = data_in[0];
			8'b00001100 : data_out[48] = data_in[0];
			8'b10001100 : data_out[49] = data_in[0];
			8'b01001100 : data_out[50] = data_in[0];
			8'b11001100 : data_out[51] = data_in[0];
			8'b00101100 : data_out[52] = data_in[0];
			8'b10101100 : data_out[53] = data_in[0];
			8'b01101100 : data_out[54] = data_in[0];
			8'b11101100 : data_out[55] = data_in[0];
			8'b00011100 : data_out[56] = data_in[0];
			8'b10011100 : data_out[57] = data_in[0];
			8'b01011100 : data_out[58] = data_in[0];
			8'b11011100 : data_out[59] = data_in[0];
			8'b00111100 : data_out[60] = data_in[0];
			8'b10111100 : data_out[61] = data_in[0];
			8'b01111100 : data_out[62] = data_in[0];
			8'b11111100 : data_out[63] = data_in[0];
			8'b00000010 : data_out[64] = data_in[0];
			8'b10000010 : data_out[65] = data_in[0];
			8'b01000010 : data_out[66] = data_in[0];
			8'b11000010 : data_out[67] = data_in[0];
			8'b00100010 : data_out[68] = data_in[0];
			8'b10100010 : data_out[69] = data_in[0];
			8'b01100010 : data_out[70] = data_in[0];
			8'b11100010 : data_out[71] = data_in[0];
			8'b00010010 : data_out[72] = data_in[0];
			8'b10010010 : data_out[73] = data_in[0];
			8'b01010010 : data_out[74] = data_in[0];
			8'b11010010 : data_out[75] = data_in[0];
			8'b00110010 : data_out[76] = data_in[0];
			8'b10110010 : data_out[77] = data_in[0];
			8'b01110010 : data_out[78] = data_in[0];
			8'b11110010 : data_out[79] = data_in[0];
			8'b00001010 : data_out[80] = data_in[0];
			8'b10001010 : data_out[81] = data_in[0];
			8'b01001010 : data_out[82] = data_in[0];
			8'b11001010 : data_out[83] = data_in[0];
			8'b00101010 : data_out[84] = data_in[0];
			8'b10101010 : data_out[85] = data_in[0];
			8'b01101010 : data_out[86] = data_in[0];
			8'b11101010 : data_out[87] = data_in[0];
			8'b00011010 : data_out[88] = data_in[0];
			8'b10011010 : data_out[89] = data_in[0];
			8'b01011010 : data_out[90] = data_in[0];
			8'b11011010 : data_out[91] = data_in[0];
			8'b00111010 : data_out[92] = data_in[0];
			8'b10111010 : data_out[93] = data_in[0];
			8'b01111010 : data_out[94] = data_in[0];
			8'b11111010 : data_out[95] = data_in[0];
			8'b00000110 : data_out[96] = data_in[0];
			8'b10000110 : data_out[97] = data_in[0];
			8'b01000110 : data_out[98] = data_in[0];
			8'b11000110 : data_out[99] = data_in[0];
			8'b00100110 : data_out[100] = data_in[0];
			8'b10100110 : data_out[101] = data_in[0];
			8'b01100110 : data_out[102] = data_in[0];
			8'b11100110 : data_out[103] = data_in[0];
			8'b00010110 : data_out[104] = data_in[0];
			8'b10010110 : data_out[105] = data_in[0];
			8'b01010110 : data_out[106] = data_in[0];
			8'b11010110 : data_out[107] = data_in[0];
			8'b00110110 : data_out[108] = data_in[0];
			8'b10110110 : data_out[109] = data_in[0];
			8'b01110110 : data_out[110] = data_in[0];
			8'b11110110 : data_out[111] = data_in[0];
			8'b00001110 : data_out[112] = data_in[0];
			8'b10001110 : data_out[113] = data_in[0];
			8'b01001110 : data_out[114] = data_in[0];
			8'b11001110 : data_out[115] = data_in[0];
			8'b00101110 : data_out[116] = data_in[0];
			8'b10101110 : data_out[117] = data_in[0];
			8'b01101110 : data_out[118] = data_in[0];
			8'b11101110 : data_out[119] = data_in[0];
			8'b00011110 : data_out[120] = data_in[0];
			8'b10011110 : data_out[121] = data_in[0];
			8'b01011110 : data_out[122] = data_in[0];
			8'b11011110 : data_out[123] = data_in[0];
			8'b00111110 : data_out[124] = data_in[0];
			8'b10111110 : data_out[125] = data_in[0];
			8'b01111110 : data_out[126] = data_in[0];
			8'b11111110 : data_out[127] = data_in[0];
			8'b00000001 : data_out[128] = data_in[0];
			8'b10000001 : data_out[129] = data_in[0];
			8'b01000001 : data_out[130] = data_in[0];
			8'b11000001 : data_out[131] = data_in[0];
			8'b00100001 : data_out[132] = data_in[0];
			8'b10100001 : data_out[133] = data_in[0];
			8'b01100001 : data_out[134] = data_in[0];
			8'b11100001 : data_out[135] = data_in[0];
			8'b00010001 : data_out[136] = data_in[0];
			8'b10010001 : data_out[137] = data_in[0];
			8'b01010001 : data_out[138] = data_in[0];
			8'b11010001 : data_out[139] = data_in[0];
			8'b00110001 : data_out[140] = data_in[0];
			8'b10110001 : data_out[141] = data_in[0];
			8'b01110001 : data_out[142] = data_in[0];
			8'b11110001 : data_out[143] = data_in[0];
			8'b00001001 : data_out[144] = data_in[0];
			8'b10001001 : data_out[145] = data_in[0];
			8'b01001001 : data_out[146] = data_in[0];
			8'b11001001 : data_out[147] = data_in[0];
			8'b00101001 : data_out[148] = data_in[0];
			8'b10101001 : data_out[149] = data_in[0];
			8'b01101001 : data_out[150] = data_in[0];
			8'b11101001 : data_out[151] = data_in[0];
			8'b00011001 : data_out[152] = data_in[0];
			8'b10011001 : data_out[153] = data_in[0];
			8'b01011001 : data_out[154] = data_in[0];
			8'b11011001 : data_out[155] = data_in[0];
			8'b00111001 : data_out[156] = data_in[0];
			8'b10111001 : data_out[157] = data_in[0];
			8'b01111001 : data_out[158] = data_in[0];
			8'b11111001 : data_out[159] = data_in[0];
			8'b00000101 : data_out[160] = data_in[0];
			8'b10000101 : data_out[161] = data_in[0];
			8'b01000101 : data_out[162] = data_in[0];
			8'b11000101 : data_out[163] = data_in[0];
			8'b00100101 : data_out[164] = data_in[0];
			8'b10100101 : data_out[165] = data_in[0];
			8'b01100101 : data_out[166] = data_in[0];
			8'b11100101 : data_out[167] = data_in[0];
			8'b00010101 : data_out[168] = data_in[0];
			8'b10010101 : data_out[169] = data_in[0];
			8'b01010101 : data_out[170] = data_in[0];
			8'b11010101 : data_out[171] = data_in[0];
			8'b00110101 : data_out[172] = data_in[0];
			8'b10110101 : data_out[173] = data_in[0];
			8'b01110101 : data_out[174] = data_in[0];
			8'b11110101 : data_out[175] = data_in[0];
			8'b00001101 : data_out[176] = data_in[0];
			8'b10001101 : data_out[177] = data_in[0];
			8'b01001101 : data_out[178] = data_in[0];
			default : 		data_out[0:178] = {179{1'bz}};
		endcase
	end
	else begin
		data_out[0:178] = {179{1'bz}};
	end
end
// ----- END Verilog codes for Decoder convert 8-bit addr to 179-bit data -----
endmodule
// ----- END Verilog module for decoder_with_data_in_8to179 -----

//----- Default net type -----
// `default_nettype none

//----- Default net type -----
// `default_nettype wire

// ----- Verilog module for decoder8to179 -----
module decoder8to179(enable,
                     address,
                     data_out);
//----- INPUT PORTS -----
input [0:0] enable;
//----- INPUT PORTS -----
input [0:7] address;
//----- OUTPUT PORTS -----
output [0:178] data_out;

//----- BEGIN Registered ports -----
reg [0:178] data_out;
//----- END Registered ports -----

// ----- BEGIN Verilog codes for Decoder convert 8-bit addr to 179-bit data -----
always@(address[0:7] or enable[0]) begin
	if (enable[0] == 1'b1) begin
		case (address[0:7])
			{8{1'b0}} : data_out[0:178] = 179'b10000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10000000 : data_out[0:178] = 179'b01000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01000000 : data_out[0:178] = 179'b00100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11000000 : data_out[0:178] = 179'b00010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00100000 : data_out[0:178] = 179'b00001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10100000 : data_out[0:178] = 179'b00000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01100000 : data_out[0:178] = 179'b00000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11100000 : data_out[0:178] = 179'b00000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00010000 : data_out[0:178] = 179'b00000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10010000 : data_out[0:178] = 179'b00000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01010000 : data_out[0:178] = 179'b00000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11010000 : data_out[0:178] = 179'b00000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00110000 : data_out[0:178] = 179'b00000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10110000 : data_out[0:178] = 179'b00000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01110000 : data_out[0:178] = 179'b00000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11110000 : data_out[0:178] = 179'b00000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00001000 : data_out[0:178] = 179'b00000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10001000 : data_out[0:178] = 179'b00000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01001000 : data_out[0:178] = 179'b00000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11001000 : data_out[0:178] = 179'b00000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00101000 : data_out[0:178] = 179'b00000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10101000 : data_out[0:178] = 179'b00000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01101000 : data_out[0:178] = 179'b00000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11101000 : data_out[0:178] = 179'b00000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00011000 : data_out[0:178] = 179'b00000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10011000 : data_out[0:178] = 179'b00000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01011000 : data_out[0:178] = 179'b00000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11011000 : data_out[0:178] = 179'b00000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00111000 : data_out[0:178] = 179'b00000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10111000 : data_out[0:178] = 179'b00000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01111000 : data_out[0:178] = 179'b00000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11111000 : data_out[0:178] = 179'b00000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00000100 : data_out[0:178] = 179'b00000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10000100 : data_out[0:178] = 179'b00000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01000100 : data_out[0:178] = 179'b00000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11000100 : data_out[0:178] = 179'b00000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00100100 : data_out[0:178] = 179'b00000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10100100 : data_out[0:178] = 179'b00000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01100100 : data_out[0:178] = 179'b00000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11100100 : data_out[0:178] = 179'b00000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00010100 : data_out[0:178] = 179'b00000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10010100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01010100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11010100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00110100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10110100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01110100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11110100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00001100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10001100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01001100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11001100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00101100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10101100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01101100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11101100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00011100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10011100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01011100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11011100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00111100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10111100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01111100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11111100 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00000010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10000010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01000010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11000010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00100010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10100010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01100010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11100010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00010010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10010010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01010010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11010010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00110010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10110010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01110010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11110010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00001010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10001010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01001010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11001010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00101010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10101010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01101010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11101010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00011010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10011010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01011010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11011010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00111010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10111010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01111010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11111010 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00000110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10000110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01000110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11000110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00100110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10100110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01100110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11100110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00010110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10010110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01010110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000;
			8'b11010110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000;
			8'b00110110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000;
			8'b10110110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000;
			8'b01110110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000;
			8'b11110110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000;
			8'b00001110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000;
			8'b10001110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000;
			8'b01001110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000;
			8'b11001110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000;
			8'b00101110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000;
			8'b10101110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000;
			8'b01101110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000;
			8'b11101110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000;
			8'b00011110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000;
			8'b10011110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000;
			8'b01011110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000;
			8'b11011110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000;
			8'b00111110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000;
			8'b10111110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000;
			8'b01111110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000;
			8'b11111110 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000;
			8'b00000001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000;
			8'b10000001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000;
			8'b01000001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000;
			8'b11000001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000;
			8'b00100001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000;
			8'b10100001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000;
			8'b01100001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000;
			8'b11100001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000;
			8'b00010001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000;
			8'b10010001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000;
			8'b01010001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000;
			8'b11010001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000;
			8'b00110001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000;
			8'b10110001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000;
			8'b01110001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000;
			8'b11110001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000;
			8'b00001001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000;
			8'b10001001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000;
			8'b01001001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000;
			8'b11001001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000;
			8'b00101001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000;
			8'b10101001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000;
			8'b01101001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000;
			8'b11101001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000;
			8'b00011001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000;
			8'b10011001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000;
			8'b01011001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000;
			8'b11011001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000;
			8'b00111001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000;
			8'b10111001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000;
			8'b01111001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000;
			8'b11111001 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000;
			8'b00000101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000;
			8'b10000101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000;
			8'b01000101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000;
			8'b11000101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000;
			8'b00100101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000;
			8'b10100101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000;
			8'b01100101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000;
			8'b11100101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000;
			8'b00010101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000;
			8'b10010101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000;
			8'b01010101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000;
			8'b11010101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000;
			8'b00110101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000;
			8'b10110101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000;
			8'b01110101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000;
			8'b11110101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000;
			8'b00001101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100;
			8'b10001101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010;
			8'b01001101 : data_out[0:178] = 179'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
			default : data_out[0:178] = {179{1'b0}};
		endcase
	end
	else begin
		data_out[0:178] = {179{1'b0}};
	end
end
// ----- END Verilog codes for Decoder convert 8-bit addr to 179-bit data -----
endmodule
// ----- END Verilog module for decoder8to179 -----

//----- Default net type -----
// `default_nettype none

