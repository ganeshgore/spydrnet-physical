//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Thu Oct 28 18:40:07 2021
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
// `default_nettype wire

// ----- Verilog module for fpga_top -----
module fpga_top(cfg_done,
                prog_reset,
                prog_clk,
                reset,
                clk,
                gfpga_pad_GPIO_PAD,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] cfg_done;
//----- GLOBAL PORTS -----
input [0:0] prog_reset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] reset;
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GPIO PORTS -----
inout [0:127] gfpga_pad_GPIO_PAD;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:19] cbx_1__0__0_chanx_left_out;
wire [0:19] cbx_1__0__0_chanx_right_out;
wire [0:19] cbx_1__0__1_chanx_left_out;
wire [0:19] cbx_1__0__1_chanx_right_out;
wire [0:19] cbx_1__0__2_chanx_left_out;
wire [0:19] cbx_1__0__2_chanx_right_out;
wire [0:19] cbx_1__0__3_chanx_left_out;
wire [0:19] cbx_1__0__3_chanx_right_out;
wire [0:19] cbx_1__1__0_chanx_left_out;
wire [0:19] cbx_1__1__0_chanx_right_out;
wire [0:19] cbx_1__1__10_chanx_left_out;
wire [0:19] cbx_1__1__10_chanx_right_out;
wire [0:19] cbx_1__1__11_chanx_left_out;
wire [0:19] cbx_1__1__11_chanx_right_out;
wire [0:19] cbx_1__1__1_chanx_left_out;
wire [0:19] cbx_1__1__1_chanx_right_out;
wire [0:19] cbx_1__1__2_chanx_left_out;
wire [0:19] cbx_1__1__2_chanx_right_out;
wire [0:19] cbx_1__1__3_chanx_left_out;
wire [0:19] cbx_1__1__3_chanx_right_out;
wire [0:19] cbx_1__1__4_chanx_left_out;
wire [0:19] cbx_1__1__4_chanx_right_out;
wire [0:19] cbx_1__1__5_chanx_left_out;
wire [0:19] cbx_1__1__5_chanx_right_out;
wire [0:19] cbx_1__1__6_chanx_left_out;
wire [0:19] cbx_1__1__6_chanx_right_out;
wire [0:19] cbx_1__1__7_chanx_left_out;
wire [0:19] cbx_1__1__7_chanx_right_out;
wire [0:19] cbx_1__1__8_chanx_left_out;
wire [0:19] cbx_1__1__8_chanx_right_out;
wire [0:19] cbx_1__1__9_chanx_left_out;
wire [0:19] cbx_1__1__9_chanx_right_out;
wire [0:19] cbx_1__4__0_chanx_left_out;
wire [0:19] cbx_1__4__0_chanx_right_out;
wire [0:19] cbx_1__4__1_chanx_left_out;
wire [0:19] cbx_1__4__1_chanx_right_out;
wire [0:19] cbx_1__4__2_chanx_left_out;
wire [0:19] cbx_1__4__2_chanx_right_out;
wire [0:19] cbx_1__4__3_chanx_left_out;
wire [0:19] cbx_1__4__3_chanx_right_out;
wire [0:19] cby_0__1__0_chany_bottom_out;
wire [0:19] cby_0__1__0_chany_top_out;
wire [0:19] cby_0__1__1_chany_bottom_out;
wire [0:19] cby_0__1__1_chany_top_out;
wire [0:19] cby_0__1__2_chany_bottom_out;
wire [0:19] cby_0__1__2_chany_top_out;
wire [0:19] cby_0__1__3_chany_bottom_out;
wire [0:19] cby_0__1__3_chany_top_out;
wire [0:19] cby_1__1__0_chany_bottom_out;
wire [0:19] cby_1__1__0_chany_top_out;
wire [0:19] cby_1__1__10_chany_bottom_out;
wire [0:19] cby_1__1__10_chany_top_out;
wire [0:19] cby_1__1__11_chany_bottom_out;
wire [0:19] cby_1__1__11_chany_top_out;
wire [0:19] cby_1__1__1_chany_bottom_out;
wire [0:19] cby_1__1__1_chany_top_out;
wire [0:19] cby_1__1__2_chany_bottom_out;
wire [0:19] cby_1__1__2_chany_top_out;
wire [0:19] cby_1__1__3_chany_bottom_out;
wire [0:19] cby_1__1__3_chany_top_out;
wire [0:19] cby_1__1__4_chany_bottom_out;
wire [0:19] cby_1__1__4_chany_top_out;
wire [0:19] cby_1__1__5_chany_bottom_out;
wire [0:19] cby_1__1__5_chany_top_out;
wire [0:19] cby_1__1__6_chany_bottom_out;
wire [0:19] cby_1__1__6_chany_top_out;
wire [0:19] cby_1__1__7_chany_bottom_out;
wire [0:19] cby_1__1__7_chany_top_out;
wire [0:19] cby_1__1__8_chany_bottom_out;
wire [0:19] cby_1__1__8_chany_top_out;
wire [0:19] cby_1__1__9_chany_bottom_out;
wire [0:19] cby_1__1__9_chany_top_out;
wire [0:19] cby_4__1__0_chany_bottom_out;
wire [0:19] cby_4__1__0_chany_top_out;
wire [0:19] cby_4__1__1_chany_bottom_out;
wire [0:19] cby_4__1__1_chany_top_out;
wire [0:19] cby_4__1__2_chany_bottom_out;
wire [0:19] cby_4__1__2_chany_top_out;
wire [0:19] cby_4__1__3_chany_bottom_out;
wire [0:19] cby_4__1__3_chany_top_out;
wire [0:19] sb_0__0__0_chanx_right_out;
wire [0:19] sb_0__0__0_chany_top_out;
wire [0:19] sb_0__1__0_chanx_right_out;
wire [0:19] sb_0__1__0_chany_bottom_out;
wire [0:19] sb_0__1__0_chany_top_out;
wire [0:19] sb_0__1__1_chanx_right_out;
wire [0:19] sb_0__1__1_chany_bottom_out;
wire [0:19] sb_0__1__1_chany_top_out;
wire [0:19] sb_0__1__2_chanx_right_out;
wire [0:19] sb_0__1__2_chany_bottom_out;
wire [0:19] sb_0__1__2_chany_top_out;
wire [0:19] sb_0__4__0_chanx_right_out;
wire [0:19] sb_0__4__0_chany_bottom_out;
wire [0:19] sb_1__0__0_chanx_left_out;
wire [0:19] sb_1__0__0_chanx_right_out;
wire [0:19] sb_1__0__0_chany_top_out;
wire [0:19] sb_1__0__1_chanx_left_out;
wire [0:19] sb_1__0__1_chanx_right_out;
wire [0:19] sb_1__0__1_chany_top_out;
wire [0:19] sb_1__0__2_chanx_left_out;
wire [0:19] sb_1__0__2_chanx_right_out;
wire [0:19] sb_1__0__2_chany_top_out;
wire [0:19] sb_1__1__0_chanx_left_out;
wire [0:19] sb_1__1__0_chanx_right_out;
wire [0:19] sb_1__1__0_chany_bottom_out;
wire [0:19] sb_1__1__0_chany_top_out;
wire [0:19] sb_1__1__1_chanx_left_out;
wire [0:19] sb_1__1__1_chanx_right_out;
wire [0:19] sb_1__1__1_chany_bottom_out;
wire [0:19] sb_1__1__1_chany_top_out;
wire [0:19] sb_1__1__2_chanx_left_out;
wire [0:19] sb_1__1__2_chanx_right_out;
wire [0:19] sb_1__1__2_chany_bottom_out;
wire [0:19] sb_1__1__2_chany_top_out;
wire [0:19] sb_1__1__3_chanx_left_out;
wire [0:19] sb_1__1__3_chanx_right_out;
wire [0:19] sb_1__1__3_chany_bottom_out;
wire [0:19] sb_1__1__3_chany_top_out;
wire [0:19] sb_1__1__4_chanx_left_out;
wire [0:19] sb_1__1__4_chanx_right_out;
wire [0:19] sb_1__1__4_chany_bottom_out;
wire [0:19] sb_1__1__4_chany_top_out;
wire [0:19] sb_1__1__5_chanx_left_out;
wire [0:19] sb_1__1__5_chanx_right_out;
wire [0:19] sb_1__1__5_chany_bottom_out;
wire [0:19] sb_1__1__5_chany_top_out;
wire [0:19] sb_1__1__6_chanx_left_out;
wire [0:19] sb_1__1__6_chanx_right_out;
wire [0:19] sb_1__1__6_chany_bottom_out;
wire [0:19] sb_1__1__6_chany_top_out;
wire [0:19] sb_1__1__7_chanx_left_out;
wire [0:19] sb_1__1__7_chanx_right_out;
wire [0:19] sb_1__1__7_chany_bottom_out;
wire [0:19] sb_1__1__7_chany_top_out;
wire [0:19] sb_1__1__8_chanx_left_out;
wire [0:19] sb_1__1__8_chanx_right_out;
wire [0:19] sb_1__1__8_chany_bottom_out;
wire [0:19] sb_1__1__8_chany_top_out;
wire [0:19] sb_1__4__0_chanx_left_out;
wire [0:19] sb_1__4__0_chanx_right_out;
wire [0:19] sb_1__4__0_chany_bottom_out;
wire [0:19] sb_1__4__1_chanx_left_out;
wire [0:19] sb_1__4__1_chanx_right_out;
wire [0:19] sb_1__4__1_chany_bottom_out;
wire [0:19] sb_1__4__2_chanx_left_out;
wire [0:19] sb_1__4__2_chanx_right_out;
wire [0:19] sb_1__4__2_chany_bottom_out;
wire [0:19] sb_4__0__0_chanx_left_out;
wire [0:19] sb_4__0__0_chany_top_out;
wire [0:19] sb_4__1__0_chanx_left_out;
wire [0:19] sb_4__1__0_chany_bottom_out;
wire [0:19] sb_4__1__0_chany_top_out;
wire [0:19] sb_4__1__1_chanx_left_out;
wire [0:19] sb_4__1__1_chany_bottom_out;
wire [0:19] sb_4__1__1_chany_top_out;
wire [0:19] sb_4__1__2_chanx_left_out;
wire [0:19] sb_4__1__2_chany_bottom_out;
wire [0:19] sb_4__1__2_chany_top_out;
wire [0:19] sb_4__4__0_chanx_left_out;
wire [0:19] sb_4__4__0_chany_bottom_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_clb grid_clb_1__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_0_ccff_tail));

	grid_clb grid_clb_1__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_1_ccff_tail));

	grid_clb grid_clb_1__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_2_ccff_tail));

	grid_clb grid_clb_1__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_1__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(ccff_tail));

	grid_clb grid_clb_2__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__1__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_4_ccff_tail));

	grid_clb grid_clb_2__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__1__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_5_ccff_tail));

	grid_clb grid_clb_2__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__1__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_6_ccff_tail));

	grid_clb grid_clb_2__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_2__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__1__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_7_ccff_tail));

	grid_clb grid_clb_3__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__1__8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_8_ccff_tail));

	grid_clb grid_clb_3__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__1__9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_9_ccff_tail));

	grid_clb grid_clb_3__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__1__10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_10_ccff_tail));

	grid_clb grid_clb_3__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_3__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_1__1__11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_11_ccff_tail));

	grid_clb grid_clb_4__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_4__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_12_ccff_tail));

	grid_clb grid_clb_4__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__2__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_4__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_13_ccff_tail));

	grid_clb grid_clb_4__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__3__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_4__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_14_ccff_tail));

	grid_clb grid_clb_4__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.reset(reset),
		.clk(clk),
		.top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.right_width_0_height_0_subtile_0__pin_I_13_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.right_width_0_height_0_subtile_0__pin_I_17_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.right_width_0_height_0_subtile_0__pin_I_21_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.right_width_0_height_0_subtile_0__pin_I_25_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.right_width_0_height_0_subtile_0__pin_I_29_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.right_width_0_height_0_subtile_0__pin_I_33_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.right_width_0_height_0_subtile_0__pin_I_37_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_width_0_height_0_subtile_0__pin_clk_0_(grid_clb_4__4__undriven_bottom_width_0_height_0_subtile_0__pin_clk_0_),
		.left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.ccff_head(cby_4__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_1_),
		.right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_5_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_3_),
		.left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_tail(grid_clb_15_ccff_tail));

	grid_io_top grid_io_top_1__5_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[0:7]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__4__0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_0_ccff_tail));

	grid_io_top grid_io_top_2__5_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[8:15]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__4__1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_1_ccff_tail));

	grid_io_top grid_io_top_3__5_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[16:23]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__4__2_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_2_ccff_tail));

	grid_io_top grid_io_top_4__5_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[24:31]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cbx_1__4__3_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_top_3_ccff_tail));

	grid_io_right grid_io_right_5__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[32:39]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_1_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_0_ccff_tail));

	grid_io_right grid_io_right_5__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[40:47]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_2_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_1_ccff_tail));

	grid_io_right grid_io_right_5__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[48:55]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_right_3_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_2_ccff_tail));

	grid_io_right grid_io_right_5__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[56:63]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_0_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_right_3_ccff_tail));

	grid_io_bottom grid_io_bottom_4__0_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[64:71]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_0_ccff_tail));

	grid_io_bottom grid_io_bottom_3__0_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[72:79]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_1_ccff_tail));

	grid_io_bottom grid_io_bottom_2__0_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[80:87]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(grid_io_bottom_3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_2_ccff_tail));

	grid_io_bottom grid_io_bottom_1__0_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[88:95]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_3_ccff_tail));

	grid_io_left grid_io_left_0__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[96:103]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_0_ccff_tail));

	grid_io_left grid_io_left_0__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[104:111]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_1_ccff_tail));

	grid_io_left grid_io_left_0__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[112:119]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__2_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_2_ccff_tail));

	grid_io_left grid_io_left_0__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.gfpga_pad_GPIO_PAD(gfpga_pad_GPIO_PAD[120:127]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_head(cby_0__1__3_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_tail(grid_io_left_3_ccff_tail));

	sb_0__0_ sb_0__0_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__0_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_1_ccff_tail),
		.chany_top_out(sb_0__0__0_chany_top_out[0:19]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:19]),
		.ccff_tail(sb_0__0__0_ccff_tail));

	sb_0__1_ sb_0__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__1_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__1__0_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_0_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_2_ccff_tail),
		.chany_top_out(sb_0__1__0_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__0_ccff_tail));

	sb_0__1_ sb_0__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__2_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__1__1_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_1_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_3_ccff_tail),
		.chany_top_out(sb_0__1__1_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__1_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__1_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__1_ccff_tail));

	sb_0__1_ sb_0__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__3_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__1__2_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_0__1__2_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_2_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(sb_0__4__0_ccff_tail),
		.chany_top_out(sb_0__1__2_chany_top_out[0:19]),
		.chanx_right_out(sb_0__1__2_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__1__2_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__1__2_ccff_tail));

	sb_0__4_ sb_0__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__4__0_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_0__1__3_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_left_3_right_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_top_0_ccff_tail),
		.chanx_right_out(sb_0__4__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_0__4__0_chany_bottom_out[0:19]),
		.ccff_tail(sb_0__4__0_ccff_tail));

	sb_1__0_ sb_1__0_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__0_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__0__1_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_3_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_io_left_0_ccff_tail),
		.chany_top_out(sb_1__0__0_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__0_ccff_tail));

	sb_1__0_ sb_2__0_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__4_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__0__2_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__1_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_2_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_0_ccff_tail),
		.chany_top_out(sb_1__0__1_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__1_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__1_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__1_ccff_tail));

	sb_1__0_ sb_3__0_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__8_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__0__3_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__2_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_1_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_4_ccff_tail),
		.chany_top_out(sb_1__0__2_chany_top_out[0:19]),
		.chanx_right_out(sb_1__0__2_chanx_right_out[0:19]),
		.chanx_left_out(sb_1__0__2_chanx_left_out[0:19]),
		.ccff_tail(sb_1__0__2_ccff_tail));

	sb_1__1_ sb_1__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__1_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__1__3_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_1__1__0_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__1__0_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_clb_5_ccff_tail),
		.chany_top_out(sb_1__1__0_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__0_ccff_tail));

	sb_1__1_ sb_1__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__2_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__1__4_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_1__1__1_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__1__1_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_clb_1_ccff_tail),
		.chany_top_out(sb_1__1__1_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__1_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__1_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__1_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__1_ccff_tail));

	sb_1__1_ sb_1__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__3_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__1__5_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_1__1__2_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__1__2_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_clb_7_ccff_tail),
		.chany_top_out(sb_1__1__2_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__2_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__2_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__2_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__2_ccff_tail));

	sb_1__1_ sb_2__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__5_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__1__6_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_1__1__4_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__1__3_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_clb_9_ccff_tail),
		.chany_top_out(sb_1__1__3_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__3_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__3_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__3_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__3_ccff_tail));

	sb_1__1_ sb_2__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__6_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__1__7_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_1__1__5_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__1__4_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_clb_2_ccff_tail),
		.chany_top_out(sb_1__1__4_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__4_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__4_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__4_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__4_ccff_tail));

	sb_1__1_ sb_2__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__7_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__1__8_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_1__1__6_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__1__5_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_clb_11_ccff_tail),
		.chany_top_out(sb_1__1__5_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__5_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__5_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__5_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__5_ccff_tail));

	sb_1__1_ sb_3__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__9_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__1__9_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_1__1__8_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__1__6_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_clb_13_ccff_tail),
		.chany_top_out(sb_1__1__6_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__6_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__6_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__6_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__6_ccff_tail));

	sb_1__1_ sb_3__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__10_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__1__10_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_1__1__9_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__1__7_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_clb_6_ccff_tail),
		.chany_top_out(sb_1__1__7_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__7_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__7_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__7_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__7_ccff_tail));

	sb_1__1_ sb_3__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__11_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_3_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_7_),
		.chanx_right_in(cbx_1__1__11_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_1__1__10_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__1__8_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_clb_15_ccff_tail),
		.chany_top_out(sb_1__1__8_chany_top_out[0:19]),
		.chanx_right_out(sb_1__1__8_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__1__8_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__1__8_chanx_left_out[0:19]),
		.ccff_tail(sb_1__1__8_ccff_tail));

	sb_1__4_ sb_1__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__4__1_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_1__1__3_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__4__0_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_0_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_io_top_1_ccff_tail),
		.chanx_right_out(sb_1__4__0_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__4__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__4__0_chanx_left_out[0:19]),
		.ccff_tail(sb_1__4__0_ccff_tail));

	sb_1__4_ sb_2__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__4__2_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_1__1__7_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__4__1_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_1_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_io_top_2_ccff_tail),
		.chanx_right_out(sb_1__4__1_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__4__1_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__4__1_chanx_left_out[0:19]),
		.ccff_tail(sb_1__4__1_ccff_tail));

	sb_1__4_ sb_3__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__4__3_chanx_left_out[0:19]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_8_),
		.chany_bottom_in(cby_1__1__11_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_3_),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_left_width_0_height_0_subtile_0__pin_O_7_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__4__2_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_2_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_io_top_3_ccff_tail),
		.chanx_right_out(sb_1__4__2_chanx_right_out[0:19]),
		.chany_bottom_out(sb_1__4__2_chany_bottom_out[0:19]),
		.chanx_left_out(sb_1__4__2_chanx_left_out[0:19]),
		.ccff_tail(sb_1__4__2_ccff_tail));

	sb_4__0_ sb_4__0_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__0_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__3_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_bottom_0_top_width_0_height_0_subtile_7__pin_inpad_0_),
		.ccff_head(grid_clb_8_ccff_tail),
		.chany_top_out(sb_4__0__0_chany_top_out[0:19]),
		.chanx_left_out(sb_4__0__0_chanx_left_out[0:19]),
		.ccff_tail(sb_4__0__0_ccff_tail));

	sb_4__1_ sb_4__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__1_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_4__1__0_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_3_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__1__9_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_clb_12_ccff_tail),
		.chany_top_out(sb_4__1__0_chany_top_out[0:19]),
		.chany_bottom_out(sb_4__1__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_4__1__0_chanx_left_out[0:19]),
		.ccff_tail(sb_4__1__0_ccff_tail));

	sb_4__1_ sb_4__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__2_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_4__1__1_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_2_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__1__10_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_clb_10_ccff_tail),
		.chany_top_out(sb_4__1__1_chany_top_out[0:19]),
		.chany_bottom_out(sb_4__1__1_chany_bottom_out[0:19]),
		.chanx_left_out(sb_4__1__1_chanx_left_out[0:19]),
		.ccff_tail(sb_4__1__1_ccff_tail));

	sb_4__1_ sb_4__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_4__1__3_chany_bottom_out[0:19]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_1_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_5_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.chany_bottom_in(cby_4__1__2_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_1_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__1__11_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_2_),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_clb_14_ccff_tail),
		.chany_top_out(sb_4__1__2_chany_top_out[0:19]),
		.chany_bottom_out(sb_4__1__2_chany_bottom_out[0:19]),
		.chanx_left_out(sb_4__1__2_chanx_left_out[0:19]),
		.ccff_tail(sb_4__1__2_ccff_tail));

	sb_4__4_ sb_4__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_4__1__3_chany_top_out[0:19]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_4__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_5__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_6__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_right_0_left_width_0_height_0_subtile_7__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_1_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_5_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_),
		.chanx_left_in(cbx_1__4__3_chanx_right_out[0:19]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_4__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_4__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_5__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_5__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_6__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_6__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_7__pin_inpad_0_(grid_io_top_3_bottom_width_0_height_0_subtile_7__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_8_),
		.ccff_head(grid_io_right_0_ccff_tail),
		.chany_bottom_out(sb_4__4__0_chany_bottom_out[0:19]),
		.chanx_left_out(sb_4__4__0_chanx_left_out[0:19]),
		.ccff_tail(sb_4__4__0_ccff_tail));

	cbx_1__0_ cbx_1__0_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__0__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__0__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__0_ccff_tail));

	cbx_1__0_ cbx_2__0_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__1_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__1_ccff_tail),
		.chanx_left_out(cbx_1__0__1_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__1_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__0__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__1_ccff_tail));

	cbx_1__0_ cbx_3__0_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__1_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__0__2_chanx_left_out[0:19]),
		.ccff_head(sb_1__0__2_ccff_tail),
		.chanx_left_out(cbx_1__0__2_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__2_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__0__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__2_ccff_tail));

	cbx_1__0_ cbx_4__0_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__2_chanx_right_out[0:19]),
		.chanx_right_in(sb_4__0__0_chanx_left_out[0:19]),
		.ccff_head(sb_4__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__3_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__0__3_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__0__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_4__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_5__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_6__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cbx_1__0__3_ccff_tail));

	cbx_1__1_ cbx_1__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__0_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__0_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__0_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__1__0_ccff_tail));

	cbx_1__1_ cbx_1__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__1_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__1_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__1_ccff_tail),
		.chanx_left_out(cbx_1__1__1_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__1_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__1_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__1__1_ccff_tail));

	cbx_1__1_ cbx_1__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__2_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__2_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__2_ccff_tail),
		.chanx_left_out(cbx_1__1__2_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__2_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__2_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__1__2_ccff_tail));

	cbx_1__1_ cbx_2__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__3_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__3_ccff_tail),
		.chanx_left_out(cbx_1__1__3_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__3_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__3_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__1__3_ccff_tail));

	cbx_1__1_ cbx_2__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__1_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__4_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__4_ccff_tail),
		.chanx_left_out(cbx_1__1__4_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__4_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__4_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__1__4_ccff_tail));

	cbx_1__1_ cbx_2__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__2_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__5_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__5_ccff_tail),
		.chanx_left_out(cbx_1__1__5_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__5_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__5_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__1__5_ccff_tail));

	cbx_1__1_ cbx_3__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__3_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__6_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__6_ccff_tail),
		.chanx_left_out(cbx_1__1__6_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__6_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__6_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__1__6_ccff_tail));

	cbx_1__1_ cbx_3__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__4_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__7_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__7_ccff_tail),
		.chanx_left_out(cbx_1__1__7_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__7_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__7_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__1__7_ccff_tail));

	cbx_1__1_ cbx_3__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__5_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__1__8_chanx_left_out[0:19]),
		.ccff_head(sb_1__1__8_ccff_tail),
		.chanx_left_out(cbx_1__1__8_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__8_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__8_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__1__8_ccff_tail));

	cbx_1__1_ cbx_4__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__6_chanx_right_out[0:19]),
		.chanx_right_in(sb_4__1__0_chanx_left_out[0:19]),
		.ccff_head(sb_4__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__9_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__9_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__9_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__1__9_ccff_tail));

	cbx_1__1_ cbx_4__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__7_chanx_right_out[0:19]),
		.chanx_right_in(sb_4__1__1_chanx_left_out[0:19]),
		.ccff_head(sb_4__1__1_ccff_tail),
		.chanx_left_out(cbx_1__1__10_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__10_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__10_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__1__10_ccff_tail));

	cbx_1__1_ cbx_4__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__8_chanx_right_out[0:19]),
		.chanx_right_in(sb_4__1__2_chanx_left_out[0:19]),
		.ccff_head(sb_4__1__2_ccff_tail),
		.chanx_left_out(cbx_1__1__11_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__1__11_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_2_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_6_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_10_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_14_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_18_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_22_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_26_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_30_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_34_),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_(cbx_1__1__11_top_grid_bottom_width_0_height_0_subtile_0__pin_I_38_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__1__11_ccff_tail));

	cbx_1__4_ cbx_1__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__4__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__4__0_chanx_left_out[0:19]),
		.ccff_head(sb_1__4__0_ccff_tail),
		.chanx_left_out(cbx_1__4__0_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__4__0_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__4__0_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__4__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__4__0_ccff_tail));

	cbx_1__4_ cbx_2__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__0_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__4__1_chanx_left_out[0:19]),
		.ccff_head(sb_1__4__1_ccff_tail),
		.chanx_left_out(cbx_1__4__1_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__4__1_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__4__1_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__4__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__4__1_ccff_tail));

	cbx_1__4_ cbx_3__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__1_chanx_right_out[0:19]),
		.chanx_right_in(sb_1__4__2_chanx_left_out[0:19]),
		.ccff_head(sb_1__4__2_ccff_tail),
		.chanx_left_out(cbx_1__4__2_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__4__2_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__4__2_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__4__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__4__2_ccff_tail));

	cbx_1__4_ cbx_4__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__4__2_chanx_right_out[0:19]),
		.chanx_right_in(sb_4__4__0_chanx_left_out[0:19]),
		.ccff_head(sb_4__4__0_ccff_tail),
		.chanx_left_out(cbx_1__4__3_chanx_left_out[0:19]),
		.chanx_right_out(cbx_1__4__3_chanx_right_out[0:19]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_4__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_5__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_6__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_(cbx_1__4__3_top_grid_bottom_width_0_height_0_subtile_7__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_4_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_8_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_12_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_16_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_20_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_24_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_28_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_32_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_(cbx_1__4__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I_36_),
		.ccff_tail(cbx_1__4__3_ccff_tail));

	cby_0__1_ cby_0__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__0__0_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:19]),
		.ccff_head(sb_0__0__0_ccff_tail),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_0__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__0_ccff_tail));

	cby_0__1_ cby_0__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__0_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__1_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__0_ccff_tail),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_0__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__1_ccff_tail));

	cby_0__1_ cby_0__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__1_chany_top_out[0:19]),
		.chany_top_in(sb_0__1__2_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__1_ccff_tail),
		.chany_bottom_out(cby_0__1__2_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__2_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_0__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__2_ccff_tail));

	cby_0__1_ cby_0__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__2_chany_top_out[0:19]),
		.chany_top_in(sb_0__4__0_chany_bottom_out[0:19]),
		.ccff_head(sb_0__1__2_ccff_tail),
		.chany_bottom_out(cby_0__1__3_chany_bottom_out[0:19]),
		.chany_top_out(cby_0__1__3_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_0__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_4__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_5__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_6__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_7__pin_outpad_0_),
		.ccff_tail(cby_0__1__3_ccff_tail));

	cby_1__1_ cby_1__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__0_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__0__0_ccff_tail),
		.chany_bottom_out(cby_1__1__0_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__0_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__0_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__1__0_ccff_tail));

	cby_1__1_ cby_1__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__0_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__1_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__1__0_ccff_tail),
		.chany_bottom_out(cby_1__1__1_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__1_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__1_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__1__1_ccff_tail));

	cby_1__1_ cby_1__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__1_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__2_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__1__1_ccff_tail),
		.chany_bottom_out(cby_1__1__2_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__2_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__2_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__1__2_ccff_tail));

	cby_1__1_ cby_1__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__2_chany_top_out[0:19]),
		.chany_top_in(sb_1__4__0_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__1__2_ccff_tail),
		.chany_bottom_out(cby_1__1__3_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__3_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__3_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__1__3_ccff_tail));

	cby_1__1_ cby_2__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__1_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__3_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__0__1_ccff_tail),
		.chany_bottom_out(cby_1__1__4_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__4_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__4_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__1__4_ccff_tail));

	cby_1__1_ cby_2__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__3_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__4_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__1__3_ccff_tail),
		.chany_bottom_out(cby_1__1__5_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__5_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__5_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__1__5_ccff_tail));

	cby_1__1_ cby_2__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__4_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__5_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__1__4_ccff_tail),
		.chany_bottom_out(cby_1__1__6_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__6_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__6_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__1__6_ccff_tail));

	cby_1__1_ cby_2__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__5_chany_top_out[0:19]),
		.chany_top_in(sb_1__4__1_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__1__5_ccff_tail),
		.chany_bottom_out(cby_1__1__7_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__7_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__7_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__1__7_ccff_tail));

	cby_1__1_ cby_3__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__2_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__6_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__0__2_ccff_tail),
		.chany_bottom_out(cby_1__1__8_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__8_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__8_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__1__8_ccff_tail));

	cby_1__1_ cby_3__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__6_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__7_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__1__6_ccff_tail),
		.chany_bottom_out(cby_1__1__9_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__9_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__9_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__1__9_ccff_tail));

	cby_1__1_ cby_3__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__7_chany_top_out[0:19]),
		.chany_top_in(sb_1__1__8_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__1__7_ccff_tail),
		.chany_bottom_out(cby_1__1__10_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__10_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__10_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__1__10_ccff_tail));

	cby_1__1_ cby_3__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__8_chany_top_out[0:19]),
		.chany_top_in(sb_1__4__2_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__1__8_ccff_tail),
		.chany_bottom_out(cby_1__1__11_chany_bottom_out[0:19]),
		.chany_top_out(cby_1__1__11_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_3_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_3_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_7_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_7_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_11_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_11_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_15_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_15_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_19_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_19_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_23_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_23_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_27_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_27_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_31_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_31_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_35_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_35_),
		.right_grid_left_width_0_height_0_subtile_0__pin_I_39_(cby_1__1__11_right_grid_left_width_0_height_0_subtile_0__pin_I_39_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_1__1__11_ccff_tail));

	cby_4__1_ cby_4__1_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__0__0_chany_top_out[0:19]),
		.chany_top_in(sb_4__1__0_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__0__3_ccff_tail),
		.chany_bottom_out(cby_4__1__0_chany_bottom_out[0:19]),
		.chany_top_out(cby_4__1__0_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__0_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_4__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_4__1__0_ccff_tail));

	cby_4__1_ cby_4__2_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__0_chany_top_out[0:19]),
		.chany_top_in(sb_4__1__1_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__1__9_ccff_tail),
		.chany_bottom_out(cby_4__1__1_chany_bottom_out[0:19]),
		.chany_top_out(cby_4__1__1_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__1_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_4__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_4__1__1_ccff_tail));

	cby_4__1_ cby_4__3_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__1_chany_top_out[0:19]),
		.chany_top_in(sb_4__1__2_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__1__10_ccff_tail),
		.chany_bottom_out(cby_4__1__2_chany_bottom_out[0:19]),
		.chany_top_out(cby_4__1__2_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__2_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_4__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_4__1__2_ccff_tail));

	cby_4__1_ cby_4__4_ (
		.cfg_done(cfg_done),
		.prog_reset(prog_reset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_4__1__2_chany_top_out[0:19]),
		.chany_top_in(sb_4__4__0_chany_bottom_out[0:19]),
		.ccff_head(cbx_1__1__11_ccff_tail),
		.chany_bottom_out(cby_4__1__3_chany_bottom_out[0:19]),
		.chany_top_out(cby_4__1__3_chany_top_out[0:19]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_4__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_5__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_6__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_(cby_4__1__3_right_grid_left_width_0_height_0_subtile_7__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_1_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_5_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_5_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_9_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_9_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_13_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_13_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_17_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_17_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_21_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_21_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_25_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_25_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_29_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_29_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_33_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_33_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I_37_(cby_4__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I_37_),
		.ccff_tail(cby_4__1__3_ccff_tail));

endmodule
// ----- END Verilog module for fpga_top -----

//----- Default net type -----
// `default_nettype none




